magic
tech ihp-sg13g2
magscale 1 2
timestamp 1770223072
<< metal1 >>
rect 1152 9848 8352 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 8352 9848
rect 1152 9784 8352 9808
rect 2667 9596 2709 9605
rect 2667 9556 2668 9596
rect 2708 9556 2709 9596
rect 2667 9547 2709 9556
rect 3051 9596 3093 9605
rect 3051 9556 3052 9596
rect 3092 9556 3093 9596
rect 3051 9547 3093 9556
rect 3907 9596 3965 9597
rect 3907 9556 3916 9596
rect 3956 9556 3965 9596
rect 3907 9555 3965 9556
rect 1411 9512 1469 9513
rect 1411 9472 1420 9512
rect 1460 9472 1469 9512
rect 1411 9471 1469 9472
rect 5059 9512 5117 9513
rect 5059 9472 5068 9512
rect 5108 9472 5117 9512
rect 5059 9471 5117 9472
rect 7843 9512 7901 9513
rect 7843 9472 7852 9512
rect 7892 9472 7901 9512
rect 7843 9471 7901 9472
rect 2275 9428 2333 9429
rect 2275 9388 2284 9428
rect 2324 9388 2333 9428
rect 2275 9387 2333 9388
rect 3715 9428 3773 9429
rect 3715 9388 3724 9428
rect 3764 9388 3773 9428
rect 3715 9387 3773 9388
rect 3915 9428 3957 9437
rect 3915 9388 3916 9428
rect 3956 9388 3957 9428
rect 3915 9379 3957 9388
rect 4003 9428 4061 9429
rect 4003 9388 4012 9428
rect 4052 9388 4061 9428
rect 4003 9387 4061 9388
rect 4779 9428 4821 9437
rect 4779 9388 4780 9428
rect 4820 9388 4821 9428
rect 4779 9379 4821 9388
rect 4875 9428 4917 9437
rect 4875 9388 4876 9428
rect 4916 9388 4917 9428
rect 4875 9379 4917 9388
rect 7459 9428 7517 9429
rect 7459 9388 7468 9428
rect 7508 9388 7517 9428
rect 7459 9387 7517 9388
rect 4675 9344 4733 9345
rect 4675 9304 4684 9344
rect 4724 9304 4733 9344
rect 4675 9303 4733 9304
rect 1227 9260 1269 9269
rect 1227 9220 1228 9260
rect 1268 9220 1269 9260
rect 1227 9211 1269 9220
rect 2083 9260 2141 9261
rect 2083 9220 2092 9260
rect 2132 9220 2141 9260
rect 2083 9219 2141 9220
rect 2371 9260 2429 9261
rect 2371 9220 2380 9260
rect 2420 9220 2429 9260
rect 2371 9219 2429 9220
rect 4491 9260 4533 9269
rect 4491 9220 4492 9260
rect 4532 9220 4533 9260
rect 4491 9211 4533 9220
rect 4579 9260 4637 9261
rect 4579 9220 4588 9260
rect 4628 9220 4637 9260
rect 4579 9219 4637 9220
rect 5259 9260 5301 9269
rect 5259 9220 5260 9260
rect 5300 9220 5301 9260
rect 5259 9211 5301 9220
rect 5739 9260 5781 9269
rect 5739 9220 5740 9260
rect 5780 9220 5781 9260
rect 5739 9211 5781 9220
rect 8043 9260 8085 9269
rect 8043 9220 8044 9260
rect 8084 9220 8085 9260
rect 8043 9211 8085 9220
rect 1152 9092 8352 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 8352 9092
rect 1152 9028 8352 9052
rect 1995 8924 2037 8933
rect 1995 8884 1996 8924
rect 2036 8884 2037 8924
rect 1995 8875 2037 8884
rect 4771 8924 4829 8925
rect 4771 8884 4780 8924
rect 4820 8884 4829 8924
rect 4771 8883 4829 8884
rect 6787 8924 6845 8925
rect 6787 8884 6796 8924
rect 6836 8884 6845 8924
rect 6787 8883 6845 8884
rect 1507 8756 1565 8757
rect 1507 8716 1516 8756
rect 1556 8716 1565 8756
rect 1507 8715 1565 8716
rect 1891 8756 1949 8757
rect 1891 8716 1900 8756
rect 1940 8716 1949 8756
rect 1891 8715 1949 8716
rect 2371 8756 2429 8757
rect 2371 8716 2380 8756
rect 2420 8716 2429 8756
rect 2371 8715 2429 8716
rect 2475 8756 2517 8765
rect 2475 8716 2476 8756
rect 2516 8716 2517 8756
rect 2475 8707 2517 8716
rect 2667 8756 2709 8765
rect 2667 8716 2668 8756
rect 2708 8716 2709 8756
rect 2667 8707 2709 8716
rect 3523 8756 3581 8757
rect 3523 8716 3532 8756
rect 3572 8716 3581 8756
rect 3523 8715 3581 8716
rect 3723 8756 3765 8765
rect 3723 8716 3724 8756
rect 3764 8716 3765 8756
rect 3723 8707 3765 8716
rect 4387 8756 4445 8757
rect 4387 8716 4396 8756
rect 4436 8716 4445 8756
rect 4387 8715 4445 8716
rect 4579 8756 4637 8757
rect 4579 8716 4588 8756
rect 4628 8716 4637 8756
rect 4579 8715 4637 8716
rect 4683 8756 4725 8765
rect 4683 8716 4684 8756
rect 4724 8716 4725 8756
rect 4683 8707 4725 8716
rect 4875 8756 4917 8765
rect 4875 8716 4876 8756
rect 4916 8716 4917 8756
rect 4875 8707 4917 8716
rect 5059 8756 5117 8757
rect 5059 8716 5068 8756
rect 5108 8716 5117 8756
rect 5059 8715 5117 8716
rect 6595 8756 6653 8757
rect 6595 8716 6604 8756
rect 6644 8716 6653 8756
rect 6595 8715 6653 8716
rect 7459 8756 7517 8757
rect 7459 8716 7468 8756
rect 7508 8716 7517 8756
rect 7459 8715 7517 8716
rect 2851 8588 2909 8589
rect 2851 8548 2860 8588
rect 2900 8548 2909 8588
rect 2851 8547 2909 8548
rect 7659 8588 7701 8597
rect 7659 8548 7660 8588
rect 7700 8548 7701 8588
rect 7659 8539 7701 8548
rect 8043 8588 8085 8597
rect 8043 8548 8044 8588
rect 8084 8548 8085 8588
rect 8043 8539 8085 8548
rect 2667 8504 2709 8513
rect 2667 8464 2668 8504
rect 2708 8464 2709 8504
rect 2667 8455 2709 8464
rect 5731 8504 5789 8505
rect 5731 8464 5740 8504
rect 5780 8464 5789 8504
rect 5731 8463 5789 8464
rect 5923 8504 5981 8505
rect 5923 8464 5932 8504
rect 5972 8464 5981 8504
rect 5923 8463 5981 8464
rect 1152 8336 8352 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 8352 8336
rect 1152 8272 8352 8296
rect 2083 7916 2141 7917
rect 2083 7876 2092 7916
rect 2132 7876 2141 7916
rect 2083 7875 2141 7876
rect 2659 7916 2717 7917
rect 2659 7876 2668 7916
rect 2708 7876 2717 7916
rect 2659 7875 2717 7876
rect 3523 7916 3581 7917
rect 3523 7876 3532 7916
rect 3572 7876 3581 7916
rect 3523 7875 3581 7876
rect 4963 7916 5021 7917
rect 4963 7876 4972 7916
rect 5012 7876 5021 7916
rect 4963 7875 5021 7876
rect 5835 7916 5877 7925
rect 5835 7876 5836 7916
rect 5876 7876 5877 7916
rect 5835 7867 5877 7876
rect 6211 7916 6269 7917
rect 6211 7876 6220 7916
rect 6260 7876 6269 7916
rect 6211 7875 6269 7876
rect 7075 7916 7133 7917
rect 7075 7876 7084 7916
rect 7124 7876 7133 7916
rect 7075 7875 7133 7876
rect 2283 7832 2325 7841
rect 2283 7792 2284 7832
rect 2324 7792 2325 7832
rect 2283 7783 2325 7792
rect 1411 7748 1469 7749
rect 1411 7708 1420 7748
rect 1460 7708 1469 7748
rect 1411 7707 1469 7708
rect 4675 7748 4733 7749
rect 4675 7708 4684 7748
rect 4724 7708 4733 7748
rect 4675 7707 4733 7708
rect 5635 7748 5693 7749
rect 5635 7708 5644 7748
rect 5684 7708 5693 7748
rect 5635 7707 5693 7708
rect 8227 7748 8285 7749
rect 8227 7708 8236 7748
rect 8276 7708 8285 7748
rect 8227 7707 8285 7708
rect 1152 7580 8352 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 8352 7580
rect 1152 7516 8352 7540
rect 5547 7454 5589 7463
rect 5547 7414 5548 7454
rect 5588 7414 5589 7454
rect 5547 7405 5589 7414
rect 8227 7412 8285 7413
rect 8227 7372 8236 7412
rect 8276 7372 8285 7412
rect 8227 7371 8285 7372
rect 2187 7328 2229 7337
rect 2187 7288 2188 7328
rect 2228 7288 2229 7328
rect 2187 7279 2229 7288
rect 5059 7328 5117 7329
rect 5059 7288 5068 7328
rect 5108 7288 5117 7328
rect 5059 7287 5117 7288
rect 5835 7328 5877 7337
rect 5835 7288 5836 7328
rect 5876 7288 5877 7328
rect 5835 7279 5877 7288
rect 2563 7244 2621 7245
rect 2563 7204 2572 7244
rect 2612 7204 2621 7244
rect 2563 7203 2621 7204
rect 3427 7244 3485 7245
rect 3427 7204 3436 7244
rect 3476 7204 3485 7244
rect 3427 7203 3485 7204
rect 5259 7244 5301 7253
rect 5259 7204 5260 7244
rect 5300 7204 5301 7244
rect 5259 7195 5301 7204
rect 5355 7244 5397 7253
rect 5355 7204 5356 7244
rect 5396 7204 5397 7244
rect 5355 7195 5397 7204
rect 6211 7244 6269 7245
rect 6211 7204 6220 7244
rect 6260 7204 6269 7244
rect 6211 7203 6269 7204
rect 7075 7244 7133 7245
rect 7075 7204 7084 7244
rect 7124 7204 7133 7244
rect 7075 7203 7133 7204
rect 1411 7160 1469 7161
rect 1411 7120 1420 7160
rect 1460 7120 1469 7160
rect 1411 7119 1469 7120
rect 1603 7160 1661 7161
rect 1603 7120 1612 7160
rect 1652 7120 1661 7160
rect 1603 7119 1661 7120
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 1227 7076 1269 7085
rect 1227 7036 1228 7076
rect 1268 7036 1269 7076
rect 1227 7027 1269 7036
rect 1803 7076 1845 7085
rect 1803 7036 1804 7076
rect 1844 7036 1845 7076
rect 1803 7027 1845 7036
rect 1152 6824 8352 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 8352 6824
rect 1152 6760 8352 6784
rect 2659 6656 2717 6657
rect 2659 6616 2668 6656
rect 2708 6616 2717 6656
rect 2659 6615 2717 6616
rect 8235 6656 8277 6665
rect 8235 6616 8236 6656
rect 8276 6616 8277 6656
rect 8235 6607 8277 6616
rect 2475 6572 2517 6581
rect 2475 6532 2476 6572
rect 2516 6532 2517 6572
rect 2475 6523 2517 6532
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 6019 6488 6077 6489
rect 6019 6448 6028 6488
rect 6068 6448 6077 6488
rect 6019 6447 6077 6448
rect 8035 6488 8093 6489
rect 8035 6448 8044 6488
rect 8084 6448 8093 6488
rect 8035 6447 8093 6448
rect 1515 6404 1557 6413
rect 1515 6364 1516 6404
rect 1556 6364 1557 6404
rect 1515 6355 1557 6364
rect 1707 6404 1749 6413
rect 1707 6364 1708 6404
rect 1748 6364 1749 6404
rect 1707 6355 1749 6364
rect 1891 6404 1949 6405
rect 1891 6364 1900 6404
rect 1940 6364 1949 6404
rect 1891 6363 1949 6364
rect 2091 6404 2133 6413
rect 2091 6364 2092 6404
rect 2132 6364 2133 6404
rect 2091 6355 2133 6364
rect 3331 6404 3389 6405
rect 3331 6364 3340 6404
rect 3380 6364 3389 6404
rect 3331 6363 3389 6364
rect 4195 6404 4253 6405
rect 4195 6364 4204 6404
rect 4244 6364 4253 6404
rect 4195 6363 4253 6364
rect 4587 6404 4629 6413
rect 4587 6364 4588 6404
rect 4628 6364 4629 6404
rect 4587 6355 4629 6364
rect 4683 6404 4725 6413
rect 4683 6364 4684 6404
rect 4724 6364 4725 6404
rect 4683 6355 4725 6364
rect 4875 6404 4917 6413
rect 4875 6364 4876 6404
rect 4916 6364 4917 6404
rect 4875 6355 4917 6364
rect 4971 6404 5013 6413
rect 4971 6364 4972 6404
rect 5012 6364 5013 6404
rect 4971 6355 5013 6364
rect 5067 6404 5109 6413
rect 5067 6364 5068 6404
rect 5108 6364 5109 6404
rect 5067 6355 5109 6364
rect 5163 6404 5205 6413
rect 5163 6364 5164 6404
rect 5204 6364 5205 6404
rect 5163 6355 5205 6364
rect 7459 6404 7517 6405
rect 7459 6364 7468 6404
rect 7508 6364 7517 6404
rect 7459 6363 7517 6364
rect 7843 6404 7901 6405
rect 7843 6364 7852 6404
rect 7892 6364 7901 6404
rect 7843 6363 7901 6364
rect 1995 6320 2037 6329
rect 1995 6280 1996 6320
rect 2036 6280 2037 6320
rect 1995 6271 2037 6280
rect 3523 6236 3581 6237
rect 3523 6196 3532 6236
rect 3572 6196 3581 6236
rect 3523 6195 3581 6196
rect 4387 6236 4445 6237
rect 4387 6196 4396 6236
rect 4436 6196 4445 6236
rect 4387 6195 4445 6196
rect 7755 6236 7797 6245
rect 7755 6196 7756 6236
rect 7796 6196 7797 6236
rect 7755 6187 7797 6196
rect 1152 6068 8352 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 8352 6068
rect 1152 6004 8352 6028
rect 2379 5816 2421 5825
rect 2379 5776 2380 5816
rect 2420 5776 2421 5816
rect 2379 5767 2421 5776
rect 1707 5732 1749 5741
rect 1707 5692 1708 5732
rect 1748 5692 1749 5732
rect 1707 5683 1749 5692
rect 1899 5732 1941 5741
rect 1899 5692 1900 5732
rect 1940 5692 1941 5732
rect 1899 5683 1941 5692
rect 1995 5732 2037 5741
rect 1995 5692 1996 5732
rect 2036 5692 2037 5732
rect 1995 5683 2037 5692
rect 2187 5732 2229 5741
rect 2187 5692 2188 5732
rect 2228 5692 2229 5732
rect 2187 5683 2229 5692
rect 2475 5732 2517 5741
rect 2475 5692 2476 5732
rect 2516 5692 2517 5732
rect 2475 5683 2517 5692
rect 3331 5732 3389 5733
rect 3331 5692 3340 5732
rect 3380 5692 3389 5732
rect 3331 5691 3389 5692
rect 3619 5732 3677 5733
rect 3619 5692 3628 5732
rect 3668 5692 3677 5732
rect 3619 5691 3677 5692
rect 3723 5732 3765 5741
rect 3723 5692 3724 5732
rect 3764 5692 3765 5732
rect 3723 5683 3765 5692
rect 3915 5732 3957 5741
rect 3915 5692 3916 5732
rect 3956 5692 3957 5732
rect 3915 5683 3957 5692
rect 4099 5732 4157 5733
rect 4099 5692 4108 5732
rect 4148 5692 4157 5732
rect 4099 5691 4157 5692
rect 4779 5732 4821 5741
rect 4779 5692 4780 5732
rect 4820 5692 4821 5732
rect 4779 5683 4821 5692
rect 5635 5732 5693 5733
rect 5635 5692 5644 5732
rect 5684 5692 5693 5732
rect 5635 5691 5693 5692
rect 6499 5732 6557 5733
rect 6499 5692 6508 5732
rect 6548 5692 6557 5732
rect 6499 5691 6557 5692
rect 7363 5732 7421 5733
rect 7363 5692 7372 5732
rect 7412 5692 7421 5732
rect 7363 5691 7421 5692
rect 8227 5732 8285 5733
rect 8227 5692 8236 5732
rect 8276 5692 8285 5732
rect 8227 5691 8285 5692
rect 1315 5648 1373 5649
rect 1315 5608 1324 5648
rect 1364 5608 1373 5648
rect 1315 5607 1373 5608
rect 1987 5564 2045 5565
rect 1987 5524 1996 5564
rect 2036 5524 2045 5564
rect 1987 5523 2045 5524
rect 1515 5480 1557 5489
rect 1515 5440 1516 5480
rect 1556 5440 1557 5480
rect 1515 5431 1557 5440
rect 2659 5480 2717 5481
rect 2659 5440 2668 5480
rect 2708 5440 2717 5480
rect 2659 5439 2717 5440
rect 3915 5480 3957 5489
rect 3915 5440 3916 5480
rect 3956 5440 3957 5480
rect 3915 5431 3957 5440
rect 4963 5480 5021 5481
rect 4963 5440 4972 5480
rect 5012 5440 5021 5480
rect 4963 5439 5021 5440
rect 5827 5480 5885 5481
rect 5827 5440 5836 5480
rect 5876 5440 5885 5480
rect 5827 5439 5885 5440
rect 6691 5480 6749 5481
rect 6691 5440 6700 5480
rect 6740 5440 6749 5480
rect 6691 5439 6749 5440
rect 7555 5480 7613 5481
rect 7555 5440 7564 5480
rect 7604 5440 7613 5480
rect 7555 5439 7613 5440
rect 1152 5312 8352 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 8352 5312
rect 1152 5248 8352 5272
rect 1227 5144 1269 5153
rect 1227 5104 1228 5144
rect 1268 5104 1269 5144
rect 1227 5095 1269 5104
rect 8227 5144 8285 5145
rect 8227 5104 8236 5144
rect 8276 5104 8285 5144
rect 8227 5103 8285 5104
rect 1707 5060 1749 5069
rect 1707 5020 1708 5060
rect 1748 5020 1749 5060
rect 1707 5011 1749 5020
rect 2091 5060 2133 5069
rect 2091 5020 2092 5060
rect 2132 5020 2133 5060
rect 2091 5011 2133 5020
rect 1315 4892 1373 4893
rect 1315 4852 1324 4892
rect 1364 4852 1373 4892
rect 1315 4851 1373 4852
rect 2283 4892 2325 4901
rect 2283 4852 2284 4892
rect 2324 4852 2325 4892
rect 2283 4843 2325 4852
rect 2659 4892 2717 4893
rect 2659 4852 2668 4892
rect 2708 4852 2717 4892
rect 2659 4851 2717 4852
rect 3523 4892 3581 4893
rect 3523 4852 3532 4892
rect 3572 4852 3581 4892
rect 3523 4851 3581 4852
rect 4963 4892 5021 4893
rect 4963 4852 4972 4892
rect 5012 4852 5021 4892
rect 4963 4851 5021 4852
rect 5835 4892 5877 4901
rect 5835 4852 5836 4892
rect 5876 4852 5877 4892
rect 5835 4843 5877 4852
rect 6211 4892 6269 4893
rect 6211 4852 6220 4892
rect 6260 4852 6269 4892
rect 6211 4851 6269 4852
rect 7075 4892 7133 4893
rect 7075 4852 7084 4892
rect 7124 4852 7133 4892
rect 7075 4851 7133 4852
rect 1227 4724 1269 4733
rect 1227 4684 1228 4724
rect 1268 4684 1269 4724
rect 1227 4675 1269 4684
rect 4675 4724 4733 4725
rect 4675 4684 4684 4724
rect 4724 4684 4733 4724
rect 4675 4683 4733 4684
rect 5635 4724 5693 4725
rect 5635 4684 5644 4724
rect 5684 4684 5693 4724
rect 5635 4683 5693 4684
rect 1152 4556 8352 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 8352 4556
rect 1152 4492 8352 4516
rect 4867 4388 4925 4389
rect 4867 4348 4876 4388
rect 4916 4348 4925 4388
rect 4867 4347 4925 4348
rect 1611 4304 1653 4313
rect 1611 4264 1612 4304
rect 1652 4264 1653 4304
rect 1611 4255 1653 4264
rect 2187 4304 2229 4313
rect 2187 4264 2188 4304
rect 2228 4264 2229 4304
rect 2187 4255 2229 4264
rect 8235 4304 8277 4313
rect 8235 4264 8236 4304
rect 8276 4264 8277 4304
rect 8235 4255 8277 4264
rect 1515 4220 1557 4229
rect 1515 4180 1516 4220
rect 1556 4180 1557 4220
rect 1515 4171 1557 4180
rect 1707 4220 1749 4229
rect 1707 4180 1708 4220
rect 1748 4180 1749 4220
rect 1707 4171 1749 4180
rect 2563 4220 2621 4221
rect 2563 4180 2572 4220
rect 2612 4180 2621 4220
rect 2563 4179 2621 4180
rect 3427 4220 3485 4221
rect 3427 4180 3436 4220
rect 3476 4180 3485 4220
rect 3427 4179 3485 4180
rect 5067 4220 5109 4229
rect 5067 4180 5068 4220
rect 5108 4180 5109 4220
rect 5067 4171 5109 4180
rect 5163 4220 5205 4229
rect 5163 4180 5164 4220
rect 5204 4180 5205 4220
rect 5163 4171 5205 4180
rect 5259 4220 5301 4229
rect 5259 4180 5260 4220
rect 5300 4180 5301 4220
rect 5259 4171 5301 4180
rect 5355 4220 5397 4229
rect 5355 4180 5356 4220
rect 5396 4180 5397 4220
rect 5355 4171 5397 4180
rect 6979 4220 7037 4221
rect 6979 4180 6988 4220
rect 7028 4180 7037 4220
rect 6979 4179 7037 4180
rect 7843 4220 7901 4221
rect 7843 4180 7852 4220
rect 7892 4180 7901 4220
rect 7843 4179 7901 4180
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 4579 3968 4637 3969
rect 4579 3928 4588 3968
rect 4628 3928 4637 3968
rect 4579 3927 4637 3928
rect 1152 3800 8352 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 8352 3800
rect 1152 3736 8352 3760
rect 1227 3632 1269 3641
rect 1227 3592 1228 3632
rect 1268 3592 1269 3632
rect 1227 3583 1269 3592
rect 4971 3632 5013 3641
rect 4971 3592 4972 3632
rect 5012 3592 5013 3632
rect 4971 3583 5013 3592
rect 5739 3632 5781 3641
rect 5739 3592 5740 3632
rect 5780 3592 5781 3632
rect 5739 3583 5781 3592
rect 2475 3548 2517 3557
rect 2475 3508 2476 3548
rect 2516 3508 2517 3548
rect 2475 3499 2517 3508
rect 4491 3548 4533 3557
rect 4491 3508 4492 3548
rect 4532 3508 4533 3548
rect 4491 3499 4533 3508
rect 7851 3548 7893 3557
rect 7851 3508 7852 3548
rect 7892 3508 7893 3548
rect 7851 3499 7893 3508
rect 1411 3464 1469 3465
rect 1411 3424 1420 3464
rect 1460 3424 1469 3464
rect 1411 3423 1469 3424
rect 1987 3464 2045 3465
rect 1987 3424 1996 3464
rect 2036 3424 2045 3464
rect 1987 3423 2045 3424
rect 2859 3464 2901 3473
rect 2859 3424 2860 3464
rect 2900 3424 2901 3464
rect 2859 3415 2901 3424
rect 2379 3380 2421 3389
rect 2379 3340 2380 3380
rect 2420 3340 2421 3380
rect 2379 3331 2421 3340
rect 2563 3380 2621 3381
rect 2563 3340 2572 3380
rect 2612 3340 2621 3380
rect 2563 3339 2621 3340
rect 2763 3380 2805 3389
rect 2763 3340 2764 3380
rect 2804 3340 2805 3380
rect 2763 3331 2805 3340
rect 2955 3380 2997 3389
rect 2955 3340 2956 3380
rect 2996 3340 2997 3380
rect 2955 3331 2997 3340
rect 3139 3380 3197 3381
rect 3139 3340 3148 3380
rect 3188 3340 3197 3380
rect 3139 3339 3197 3340
rect 3819 3380 3861 3389
rect 3819 3340 3820 3380
rect 3860 3340 3861 3380
rect 3819 3331 3861 3340
rect 4011 3380 4053 3389
rect 4011 3340 4012 3380
rect 4052 3340 4053 3380
rect 4011 3331 4053 3340
rect 4107 3380 4149 3389
rect 4107 3340 4108 3380
rect 4148 3340 4149 3380
rect 4107 3331 4149 3340
rect 4203 3380 4245 3389
rect 4203 3340 4204 3380
rect 4244 3340 4245 3380
rect 4203 3331 4245 3340
rect 4299 3380 4341 3389
rect 4299 3340 4300 3380
rect 4340 3340 4341 3380
rect 4299 3331 4341 3340
rect 4483 3380 4541 3381
rect 4483 3340 4492 3380
rect 4532 3340 4541 3380
rect 4483 3339 4541 3340
rect 4683 3380 4725 3389
rect 4683 3340 4684 3380
rect 4724 3340 4725 3380
rect 4683 3331 4725 3340
rect 4771 3380 4829 3381
rect 4771 3340 4780 3380
rect 4820 3340 4829 3380
rect 4771 3339 4829 3340
rect 4971 3380 5013 3389
rect 4971 3340 4972 3380
rect 5012 3340 5013 3380
rect 4971 3331 5013 3340
rect 5163 3380 5205 3389
rect 5163 3340 5164 3380
rect 5204 3340 5205 3380
rect 5163 3331 5205 3340
rect 5251 3380 5309 3381
rect 5251 3340 5260 3380
rect 5300 3340 5309 3380
rect 5251 3339 5309 3340
rect 7459 3380 7517 3381
rect 7459 3340 7468 3380
rect 7508 3340 7517 3380
rect 7459 3339 7517 3340
rect 2187 3212 2229 3221
rect 2187 3172 2188 3212
rect 2228 3172 2229 3212
rect 2187 3163 2229 3172
rect 1152 3044 8352 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 8352 3044
rect 1152 2980 8352 3004
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 2668 9556 2708 9596
rect 3052 9556 3092 9596
rect 3916 9556 3956 9596
rect 1420 9472 1460 9512
rect 5068 9472 5108 9512
rect 7852 9472 7892 9512
rect 2284 9388 2324 9428
rect 3724 9388 3764 9428
rect 3916 9388 3956 9428
rect 4012 9388 4052 9428
rect 4780 9388 4820 9428
rect 4876 9388 4916 9428
rect 7468 9388 7508 9428
rect 4684 9304 4724 9344
rect 1228 9220 1268 9260
rect 2092 9220 2132 9260
rect 2380 9220 2420 9260
rect 4492 9220 4532 9260
rect 4588 9220 4628 9260
rect 5260 9220 5300 9260
rect 5740 9220 5780 9260
rect 8044 9220 8084 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 1996 8884 2036 8924
rect 4780 8884 4820 8924
rect 6796 8884 6836 8924
rect 1516 8716 1556 8756
rect 1900 8716 1940 8756
rect 2380 8716 2420 8756
rect 2476 8716 2516 8756
rect 2668 8716 2708 8756
rect 3532 8716 3572 8756
rect 3724 8716 3764 8756
rect 4396 8716 4436 8756
rect 4588 8716 4628 8756
rect 4684 8716 4724 8756
rect 4876 8716 4916 8756
rect 5068 8716 5108 8756
rect 6604 8716 6644 8756
rect 7468 8716 7508 8756
rect 2860 8548 2900 8588
rect 7660 8548 7700 8588
rect 8044 8548 8084 8588
rect 2668 8464 2708 8504
rect 5740 8464 5780 8504
rect 5932 8464 5972 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 2092 7876 2132 7916
rect 2668 7876 2708 7916
rect 3532 7876 3572 7916
rect 4972 7876 5012 7916
rect 5836 7876 5876 7916
rect 6220 7876 6260 7916
rect 7084 7876 7124 7916
rect 2284 7792 2324 7832
rect 1420 7708 1460 7748
rect 4684 7708 4724 7748
rect 5644 7708 5684 7748
rect 8236 7708 8276 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5548 7414 5588 7454
rect 8236 7372 8276 7412
rect 2188 7288 2228 7328
rect 5068 7288 5108 7328
rect 5836 7288 5876 7328
rect 2572 7204 2612 7244
rect 3436 7204 3476 7244
rect 5260 7204 5300 7244
rect 5356 7204 5396 7244
rect 6220 7204 6260 7244
rect 7084 7204 7124 7244
rect 1420 7120 1460 7160
rect 1612 7120 1652 7160
rect 4588 7120 4628 7160
rect 1228 7036 1268 7076
rect 1804 7036 1844 7076
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 2668 6616 2708 6656
rect 8236 6616 8276 6656
rect 2476 6532 2516 6572
rect 1612 6448 1652 6488
rect 6028 6448 6068 6488
rect 8044 6448 8084 6488
rect 1516 6364 1556 6404
rect 1708 6364 1748 6404
rect 1900 6364 1940 6404
rect 2092 6364 2132 6404
rect 3340 6364 3380 6404
rect 4204 6364 4244 6404
rect 4588 6364 4628 6404
rect 4684 6364 4724 6404
rect 4876 6364 4916 6404
rect 4972 6364 5012 6404
rect 5068 6364 5108 6404
rect 5164 6364 5204 6404
rect 7468 6364 7508 6404
rect 7852 6364 7892 6404
rect 1996 6280 2036 6320
rect 3532 6196 3572 6236
rect 4396 6196 4436 6236
rect 7756 6196 7796 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 2380 5776 2420 5816
rect 1708 5692 1748 5732
rect 1900 5692 1940 5732
rect 1996 5692 2036 5732
rect 2188 5692 2228 5732
rect 2476 5692 2516 5732
rect 3340 5692 3380 5732
rect 3628 5692 3668 5732
rect 3724 5692 3764 5732
rect 3916 5692 3956 5732
rect 4108 5692 4148 5732
rect 4780 5692 4820 5732
rect 5644 5692 5684 5732
rect 6508 5692 6548 5732
rect 7372 5692 7412 5732
rect 8236 5692 8276 5732
rect 1324 5608 1364 5648
rect 1996 5524 2036 5564
rect 1516 5440 1556 5480
rect 2668 5440 2708 5480
rect 3916 5440 3956 5480
rect 4972 5440 5012 5480
rect 5836 5440 5876 5480
rect 6700 5440 6740 5480
rect 7564 5440 7604 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 1228 5104 1268 5144
rect 8236 5104 8276 5144
rect 1708 5020 1748 5060
rect 2092 5020 2132 5060
rect 1324 4852 1364 4892
rect 2284 4852 2324 4892
rect 2668 4852 2708 4892
rect 3532 4852 3572 4892
rect 4972 4852 5012 4892
rect 5836 4852 5876 4892
rect 6220 4852 6260 4892
rect 7084 4852 7124 4892
rect 1228 4684 1268 4724
rect 4684 4684 4724 4724
rect 5644 4684 5684 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4876 4348 4916 4388
rect 1612 4264 1652 4304
rect 2188 4264 2228 4304
rect 8236 4264 8276 4304
rect 1516 4180 1556 4220
rect 1708 4180 1748 4220
rect 2572 4180 2612 4220
rect 3436 4180 3476 4220
rect 5068 4180 5108 4220
rect 5164 4180 5204 4220
rect 5260 4180 5300 4220
rect 5356 4180 5396 4220
rect 6988 4180 7028 4220
rect 7852 4180 7892 4220
rect 5836 4096 5876 4136
rect 4588 3928 4628 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1228 3592 1268 3632
rect 4972 3592 5012 3632
rect 5740 3592 5780 3632
rect 2476 3508 2516 3548
rect 4492 3508 4532 3548
rect 7852 3508 7892 3548
rect 1420 3424 1460 3464
rect 1996 3424 2036 3464
rect 2860 3424 2900 3464
rect 2380 3340 2420 3380
rect 2572 3340 2612 3380
rect 2764 3340 2804 3380
rect 2956 3340 2996 3380
rect 3148 3340 3188 3380
rect 3820 3340 3860 3380
rect 4012 3340 4052 3380
rect 4108 3340 4148 3380
rect 4204 3340 4244 3380
rect 4300 3340 4340 3380
rect 4492 3340 4532 3380
rect 4684 3340 4724 3380
rect 4780 3340 4820 3380
rect 4972 3340 5012 3380
rect 5164 3340 5204 3380
rect 5260 3340 5300 3380
rect 7468 3340 7508 3380
rect 2188 3172 2228 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal2 >>
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 2668 9596 2708 9605
rect 2572 9556 2668 9596
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 2475 9512 2517 9521
rect 2475 9472 2476 9512
rect 2516 9472 2517 9512
rect 2475 9463 2517 9472
rect 1420 9378 1460 9463
rect 2284 9428 2324 9437
rect 1996 9388 2284 9428
rect 1228 9260 1268 9269
rect 1228 8009 1268 9220
rect 1803 9260 1845 9269
rect 1803 9220 1804 9260
rect 1844 9220 1845 9260
rect 1803 9211 1845 9220
rect 1516 8756 1556 8765
rect 1516 8597 1556 8716
rect 1515 8588 1557 8597
rect 1515 8548 1516 8588
rect 1556 8548 1557 8588
rect 1515 8539 1557 8548
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1227 7832 1269 7841
rect 1227 7792 1228 7832
rect 1268 7792 1269 7832
rect 1227 7783 1269 7792
rect 1228 7076 1268 7783
rect 1420 7748 1460 7757
rect 1460 7708 1556 7748
rect 1420 7699 1460 7708
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 1228 7027 1268 7036
rect 1420 7026 1460 7111
rect 1516 6404 1556 7708
rect 1611 7664 1653 7673
rect 1611 7624 1612 7664
rect 1652 7624 1653 7664
rect 1611 7615 1653 7624
rect 1612 7160 1652 7615
rect 1612 7111 1652 7120
rect 1804 7076 1844 9211
rect 1996 8924 2036 9388
rect 2284 9379 2324 9388
rect 1996 8875 2036 8884
rect 2092 9260 2132 9269
rect 1899 8756 1941 8765
rect 1899 8716 1900 8756
rect 1940 8716 1941 8756
rect 1899 8707 1941 8716
rect 1900 7160 1940 8707
rect 2092 8252 2132 9220
rect 2379 9260 2421 9269
rect 2379 9220 2380 9260
rect 2420 9220 2421 9260
rect 2379 9211 2421 9220
rect 2380 9126 2420 9211
rect 2476 8933 2516 9463
rect 2475 8924 2517 8933
rect 2475 8884 2476 8924
rect 2516 8884 2517 8924
rect 2475 8875 2517 8884
rect 2379 8756 2421 8765
rect 2379 8716 2380 8756
rect 2420 8716 2421 8756
rect 2379 8707 2421 8716
rect 2476 8756 2516 8875
rect 2476 8707 2516 8716
rect 2380 8622 2420 8707
rect 2092 8212 2228 8252
rect 2091 8084 2133 8093
rect 2091 8044 2092 8084
rect 2132 8044 2133 8084
rect 2091 8035 2133 8044
rect 2092 7916 2132 8035
rect 2092 7867 2132 7876
rect 2188 7328 2228 8212
rect 2284 7832 2324 7841
rect 2324 7792 2516 7832
rect 2284 7783 2324 7792
rect 2188 7279 2228 7288
rect 1900 7120 2228 7160
rect 1804 6749 1844 7036
rect 1803 6740 1845 6749
rect 1803 6700 1804 6740
rect 1844 6700 1845 6740
rect 1803 6691 1845 6700
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 1516 6355 1556 6364
rect 1612 6354 1652 6439
rect 1708 6404 1748 6415
rect 1708 6329 1748 6364
rect 1804 6404 1844 6691
rect 1900 6404 1940 6413
rect 1804 6364 1900 6404
rect 1707 6320 1749 6329
rect 1707 6280 1708 6320
rect 1748 6280 1749 6320
rect 1707 6271 1749 6280
rect 1227 5732 1269 5741
rect 1227 5692 1228 5732
rect 1268 5692 1269 5732
rect 1227 5683 1269 5692
rect 1707 5732 1749 5741
rect 1707 5692 1708 5732
rect 1748 5692 1749 5732
rect 1707 5683 1749 5692
rect 1228 5144 1268 5683
rect 1324 5648 1364 5657
rect 1364 5608 1460 5648
rect 1324 5599 1364 5608
rect 1228 5095 1268 5104
rect 1323 4976 1365 4985
rect 1323 4936 1324 4976
rect 1364 4936 1365 4976
rect 1323 4927 1365 4936
rect 1324 4892 1364 4927
rect 1420 4901 1460 5608
rect 1708 5598 1748 5683
rect 1516 5480 1556 5489
rect 1556 5440 1652 5480
rect 1516 5431 1556 5440
rect 1324 4841 1364 4852
rect 1419 4892 1461 4901
rect 1419 4852 1420 4892
rect 1460 4852 1461 4892
rect 1419 4843 1461 4852
rect 1228 4724 1268 4733
rect 1268 4684 1556 4724
rect 1228 4675 1268 4684
rect 1227 4556 1269 4565
rect 1227 4516 1228 4556
rect 1268 4516 1269 4556
rect 1227 4507 1269 4516
rect 1228 3632 1268 4507
rect 1516 4220 1556 4684
rect 1612 4649 1652 5440
rect 1707 5060 1749 5069
rect 1707 5020 1708 5060
rect 1748 5020 1749 5060
rect 1707 5011 1749 5020
rect 1708 4926 1748 5011
rect 1804 4985 1844 6364
rect 1900 6355 1940 6364
rect 1996 6329 2036 6414
rect 2091 6404 2133 6413
rect 2091 6364 2092 6404
rect 2132 6364 2133 6404
rect 2091 6355 2133 6364
rect 1995 6320 2037 6329
rect 1995 6280 1996 6320
rect 2036 6280 2037 6320
rect 1995 6271 2037 6280
rect 2092 6270 2132 6355
rect 1899 6236 1941 6245
rect 1899 6196 1900 6236
rect 1940 6196 1941 6236
rect 1899 6187 1941 6196
rect 1900 5732 1940 6187
rect 2188 6152 2228 7120
rect 2476 6992 2516 7792
rect 2572 7244 2612 9556
rect 2668 9547 2708 9556
rect 3052 9596 3092 9605
rect 2668 8765 2708 8850
rect 2667 8756 2709 8765
rect 3052 8756 3092 9556
rect 3916 9596 3956 9605
rect 3956 9556 4148 9596
rect 3916 9547 3956 9556
rect 3724 9428 3764 9437
rect 3724 8933 3764 9388
rect 3916 9428 3956 9437
rect 3916 9353 3956 9388
rect 4011 9428 4053 9437
rect 4011 9388 4012 9428
rect 4052 9388 4053 9428
rect 4011 9379 4053 9388
rect 3915 9344 3957 9353
rect 3915 9304 3916 9344
rect 3956 9304 3957 9344
rect 3915 9295 3957 9304
rect 3531 8924 3573 8933
rect 3531 8884 3532 8924
rect 3572 8884 3573 8924
rect 3531 8875 3573 8884
rect 3723 8924 3765 8933
rect 3723 8884 3724 8924
rect 3764 8884 3765 8924
rect 3723 8875 3765 8884
rect 2667 8716 2668 8756
rect 2708 8716 2709 8756
rect 2667 8707 2709 8716
rect 2764 8716 3092 8756
rect 3532 8756 3572 8875
rect 3916 8765 3956 9295
rect 4012 8849 4052 9379
rect 4011 8840 4053 8849
rect 4011 8800 4012 8840
rect 4052 8800 4053 8840
rect 4011 8791 4053 8800
rect 2668 8504 2708 8513
rect 2668 8093 2708 8464
rect 2667 8084 2709 8093
rect 2667 8044 2668 8084
rect 2708 8044 2709 8084
rect 2667 8035 2709 8044
rect 2668 7916 2708 7925
rect 2764 7916 2804 8716
rect 3532 8707 3572 8716
rect 3723 8756 3765 8765
rect 3723 8716 3724 8756
rect 3764 8716 3765 8756
rect 3723 8707 3765 8716
rect 3915 8756 3957 8765
rect 3915 8716 3916 8756
rect 3956 8716 3957 8756
rect 3915 8707 3957 8716
rect 3724 8622 3764 8707
rect 2859 8588 2901 8597
rect 2859 8548 2860 8588
rect 2900 8548 2901 8588
rect 2859 8539 2901 8548
rect 3531 8588 3573 8597
rect 3531 8548 3532 8588
rect 3572 8548 3573 8588
rect 3531 8539 3573 8548
rect 2860 8454 2900 8539
rect 3532 7916 3572 8539
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 2708 7876 2804 7916
rect 3436 7876 3532 7916
rect 2668 7867 2708 7876
rect 2572 7195 2612 7204
rect 3436 7244 3476 7876
rect 3532 7867 3572 7876
rect 3436 7195 3476 7204
rect 2476 6952 2708 6992
rect 2668 6656 2708 6952
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 2668 6607 2708 6616
rect 2476 6572 2516 6581
rect 2476 6161 2516 6532
rect 3339 6488 3381 6497
rect 3339 6448 3340 6488
rect 3380 6448 3381 6488
rect 3339 6439 3381 6448
rect 3340 6404 3380 6439
rect 4108 6413 4148 9556
rect 5068 9512 5108 9521
rect 7852 9512 7892 9521
rect 5108 9472 5396 9512
rect 5068 9463 5108 9472
rect 4780 9428 4820 9437
rect 4683 9344 4725 9353
rect 4683 9304 4684 9344
rect 4724 9304 4725 9344
rect 4683 9295 4725 9304
rect 4492 9260 4532 9269
rect 4492 8924 4532 9220
rect 4588 9260 4628 9269
rect 4588 8933 4628 9220
rect 4684 9210 4724 9295
rect 4780 9185 4820 9388
rect 4875 9428 4917 9437
rect 4875 9388 4876 9428
rect 4916 9388 4917 9428
rect 4875 9379 4917 9388
rect 4876 9294 4916 9379
rect 5260 9269 5300 9354
rect 5259 9260 5301 9269
rect 5259 9220 5260 9260
rect 5300 9220 5301 9260
rect 5259 9211 5301 9220
rect 4779 9176 4821 9185
rect 4779 9136 4780 9176
rect 4820 9136 4821 9176
rect 4779 9127 4821 9136
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4780 8933 4820 9018
rect 4300 8884 4532 8924
rect 4300 7589 4340 8884
rect 4396 8756 4436 8765
rect 4492 8756 4532 8884
rect 4587 8924 4629 8933
rect 4587 8884 4588 8924
rect 4628 8884 4629 8924
rect 4587 8875 4629 8884
rect 4779 8924 4821 8933
rect 4779 8884 4780 8924
rect 4820 8884 4821 8924
rect 4779 8875 4821 8884
rect 4588 8756 4628 8765
rect 4492 8716 4588 8756
rect 4299 7580 4341 7589
rect 4299 7540 4300 7580
rect 4340 7540 4341 7580
rect 4299 7531 4341 7540
rect 4396 7505 4436 8716
rect 4588 8707 4628 8716
rect 4683 8756 4725 8765
rect 4876 8756 4916 8765
rect 4683 8716 4684 8756
rect 4724 8716 4725 8756
rect 4683 8707 4725 8716
rect 4780 8716 4876 8756
rect 4684 8622 4724 8707
rect 4491 8000 4533 8009
rect 4780 8000 4820 8716
rect 4876 8707 4916 8716
rect 5068 8756 5108 8765
rect 5068 8009 5108 8716
rect 5356 8429 5396 9472
rect 7468 9428 7508 9437
rect 7276 9388 7468 9428
rect 5740 9260 5780 9269
rect 5740 8681 5780 9220
rect 6795 9176 6837 9185
rect 6795 9136 6796 9176
rect 6836 9136 6837 9176
rect 6795 9127 6837 9136
rect 6603 8924 6645 8933
rect 6603 8884 6604 8924
rect 6644 8884 6645 8924
rect 6603 8875 6645 8884
rect 6796 8924 6836 9127
rect 6796 8875 6836 8884
rect 6604 8756 6644 8875
rect 6604 8707 6644 8716
rect 5739 8672 5781 8681
rect 5739 8632 5740 8672
rect 5780 8632 5781 8672
rect 5739 8623 5781 8632
rect 7083 8588 7125 8597
rect 7083 8548 7084 8588
rect 7124 8548 7125 8588
rect 7083 8539 7125 8548
rect 5740 8504 5780 8513
rect 5452 8464 5740 8504
rect 5355 8420 5397 8429
rect 5355 8380 5356 8420
rect 5396 8380 5397 8420
rect 5355 8371 5397 8380
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4588 7960 4820 8000
rect 5067 8000 5109 8009
rect 5067 7960 5068 8000
rect 5108 7960 5109 8000
rect 4395 7496 4437 7505
rect 4395 7456 4396 7496
rect 4436 7456 4437 7496
rect 4395 7447 4437 7456
rect 4492 7220 4532 7951
rect 4588 7328 4628 7960
rect 5067 7951 5109 7960
rect 4972 7916 5012 7925
rect 4780 7876 4972 7916
rect 4684 7748 4724 7757
rect 4684 7505 4724 7708
rect 4683 7496 4725 7505
rect 4683 7456 4684 7496
rect 4724 7456 4725 7496
rect 4683 7447 4725 7456
rect 4780 7412 4820 7876
rect 4972 7867 5012 7876
rect 5452 7748 5492 8464
rect 5740 8455 5780 8464
rect 5932 8504 5972 8513
rect 5836 7916 5876 7925
rect 5932 7916 5972 8464
rect 6507 8420 6549 8429
rect 6507 8380 6508 8420
rect 6548 8380 6549 8420
rect 6507 8371 6549 8380
rect 5876 7876 5972 7916
rect 6219 7916 6261 7925
rect 6219 7876 6220 7916
rect 6260 7876 6261 7916
rect 5836 7867 5876 7876
rect 6219 7867 6261 7876
rect 6220 7782 6260 7867
rect 5356 7708 5492 7748
rect 5644 7748 5684 7757
rect 5684 7708 5876 7748
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5163 7412 5205 7421
rect 4780 7372 5108 7412
rect 5068 7328 5108 7372
rect 5163 7372 5164 7412
rect 5204 7372 5205 7412
rect 5163 7363 5205 7372
rect 4588 7288 4916 7328
rect 4396 7180 4532 7220
rect 3340 6353 3380 6364
rect 4107 6404 4149 6413
rect 4107 6364 4108 6404
rect 4148 6364 4149 6404
rect 4107 6355 4149 6364
rect 4204 6404 4244 6413
rect 3531 6236 3573 6245
rect 3531 6196 3532 6236
rect 3572 6196 3573 6236
rect 3531 6187 3573 6196
rect 1996 6112 2228 6152
rect 2475 6152 2517 6161
rect 2475 6112 2476 6152
rect 2516 6112 2517 6152
rect 1996 5741 2036 6112
rect 2475 6103 2517 6112
rect 3532 6102 3572 6187
rect 2379 5816 2421 5825
rect 2379 5776 2380 5816
rect 2420 5776 2421 5816
rect 2379 5767 2421 5776
rect 1900 5683 1940 5692
rect 1995 5732 2037 5741
rect 1995 5692 1996 5732
rect 2036 5692 2037 5732
rect 1995 5683 2037 5692
rect 2188 5732 2228 5741
rect 1995 5564 2037 5573
rect 1995 5524 1996 5564
rect 2036 5524 2037 5564
rect 1995 5515 2037 5524
rect 1996 5430 2036 5515
rect 2092 5060 2132 5069
rect 1803 4976 1845 4985
rect 1803 4936 1804 4976
rect 1844 4936 1845 4976
rect 1803 4927 1845 4936
rect 1611 4640 1653 4649
rect 1611 4600 1612 4640
rect 1652 4600 1653 4640
rect 1611 4591 1653 4600
rect 1611 4304 1653 4313
rect 1611 4264 1612 4304
rect 1652 4264 1653 4304
rect 1804 4304 1844 4927
rect 1804 4264 1940 4304
rect 1611 4255 1653 4264
rect 1516 4171 1556 4180
rect 1612 4170 1652 4255
rect 1708 4220 1748 4229
rect 1228 3583 1268 3592
rect 1419 3464 1461 3473
rect 1419 3424 1420 3464
rect 1460 3424 1461 3464
rect 1419 3415 1461 3424
rect 1420 3330 1460 3415
rect 1708 3389 1748 4180
rect 1707 3380 1749 3389
rect 1707 3340 1708 3380
rect 1748 3340 1749 3380
rect 1707 3331 1749 3340
rect 1900 3305 1940 4264
rect 2092 4229 2132 5020
rect 2188 4724 2228 5692
rect 2380 5682 2420 5767
rect 2476 5741 2516 5826
rect 4204 5825 4244 6364
rect 4396 6236 4436 7180
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 4588 7026 4628 7111
rect 4683 7076 4725 7085
rect 4683 7036 4684 7076
rect 4724 7036 4725 7076
rect 4683 7027 4725 7036
rect 4587 6404 4629 6413
rect 4587 6364 4588 6404
rect 4628 6364 4629 6404
rect 4587 6355 4629 6364
rect 4684 6404 4724 7027
rect 4684 6355 4724 6364
rect 4876 6404 4916 7288
rect 5068 7279 5108 7288
rect 5164 7244 5204 7363
rect 5260 7244 5300 7272
rect 5164 7220 5260 7244
rect 5068 7204 5260 7220
rect 5068 7180 5204 7204
rect 5260 7195 5300 7204
rect 5356 7244 5396 7708
rect 5644 7699 5684 7708
rect 5356 7195 5396 7204
rect 5548 7454 5588 7463
rect 4971 6488 5013 6497
rect 4971 6448 4972 6488
rect 5012 6448 5013 6488
rect 4971 6439 5013 6448
rect 4876 6355 4916 6364
rect 4972 6404 5012 6439
rect 4588 6270 4628 6355
rect 4972 6353 5012 6364
rect 5068 6404 5108 7180
rect 5548 6497 5588 7414
rect 5836 7328 5876 7708
rect 5836 7279 5876 7288
rect 6220 7253 6260 7338
rect 6219 7244 6261 7253
rect 6219 7204 6220 7244
rect 6260 7204 6261 7244
rect 6219 7195 6261 7204
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 5068 6355 5108 6364
rect 5163 6404 5205 6413
rect 5163 6364 5164 6404
rect 5204 6364 5205 6404
rect 5163 6355 5205 6364
rect 5164 6270 5204 6355
rect 6028 6354 6068 6439
rect 4396 6187 4436 6196
rect 6219 6152 6261 6161
rect 6219 6112 6220 6152
rect 6260 6112 6261 6152
rect 6219 6103 6261 6112
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4203 5816 4245 5825
rect 4203 5776 4204 5816
rect 4244 5776 4245 5816
rect 4203 5767 4245 5776
rect 2475 5732 2517 5741
rect 2475 5692 2476 5732
rect 2516 5692 2517 5732
rect 2475 5683 2517 5692
rect 3340 5732 3380 5741
rect 3628 5732 3668 5741
rect 3340 5573 3380 5692
rect 3532 5692 3628 5732
rect 3339 5564 3381 5573
rect 3339 5524 3340 5564
rect 3380 5524 3381 5564
rect 3339 5515 3381 5524
rect 2668 5480 2708 5489
rect 2572 5440 2668 5480
rect 2284 4892 2324 4901
rect 2572 4892 2612 5440
rect 2668 5431 2708 5440
rect 3532 5144 3572 5692
rect 3628 5683 3668 5692
rect 3724 5732 3764 5741
rect 3724 5573 3764 5692
rect 3916 5732 3956 5741
rect 4108 5732 4148 5741
rect 3956 5692 4052 5732
rect 3916 5683 3956 5692
rect 3723 5564 3765 5573
rect 3723 5524 3724 5564
rect 3764 5524 3765 5564
rect 3723 5515 3765 5524
rect 3916 5489 3956 5574
rect 3915 5480 3957 5489
rect 3915 5440 3916 5480
rect 3956 5440 3957 5480
rect 4012 5480 4052 5692
rect 4108 5564 4148 5692
rect 4779 5732 4821 5741
rect 5644 5732 5684 5741
rect 4779 5692 4780 5732
rect 4820 5692 4821 5732
rect 4779 5683 4821 5692
rect 5452 5692 5644 5732
rect 4587 5648 4629 5657
rect 4587 5608 4588 5648
rect 4628 5608 4629 5648
rect 4587 5599 4629 5608
rect 4299 5564 4341 5573
rect 4108 5524 4244 5564
rect 4012 5440 4148 5480
rect 3915 5431 3957 5440
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3532 5104 3668 5144
rect 2667 5060 2709 5069
rect 2667 5020 2668 5060
rect 2708 5020 2709 5060
rect 2667 5011 2709 5020
rect 2955 5060 2997 5069
rect 2955 5020 2956 5060
rect 2996 5020 2997 5060
rect 2955 5011 2997 5020
rect 2324 4852 2612 4892
rect 2668 4892 2708 5011
rect 2284 4843 2324 4852
rect 2668 4843 2708 4852
rect 2763 4892 2805 4901
rect 2763 4852 2764 4892
rect 2804 4852 2805 4892
rect 2763 4843 2805 4852
rect 2188 4684 2420 4724
rect 2187 4304 2229 4313
rect 2187 4264 2188 4304
rect 2228 4264 2229 4304
rect 2187 4255 2229 4264
rect 2091 4220 2133 4229
rect 2091 4180 2092 4220
rect 2132 4180 2133 4220
rect 2091 4171 2133 4180
rect 2188 4170 2228 4255
rect 1995 4052 2037 4061
rect 1995 4012 1996 4052
rect 2036 4012 2037 4052
rect 1995 4003 2037 4012
rect 1996 3464 2036 4003
rect 2380 3557 2420 4684
rect 2571 4220 2613 4229
rect 2571 4180 2572 4220
rect 2612 4180 2613 4220
rect 2571 4171 2613 4180
rect 2572 4086 2612 4171
rect 2764 3632 2804 4843
rect 2764 3592 2900 3632
rect 2379 3548 2421 3557
rect 2379 3508 2380 3548
rect 2420 3508 2421 3548
rect 2379 3499 2421 3508
rect 2476 3548 2516 3557
rect 2516 3508 2804 3548
rect 2476 3499 2516 3508
rect 1996 3415 2036 3424
rect 2380 3380 2420 3499
rect 2380 3331 2420 3340
rect 2572 3380 2612 3391
rect 2572 3305 2612 3340
rect 2764 3380 2804 3508
rect 2860 3464 2900 3592
rect 2860 3415 2900 3424
rect 2764 3331 2804 3340
rect 2956 3380 2996 5011
rect 3532 4892 3572 4901
rect 3436 4220 3476 4229
rect 3532 4220 3572 4852
rect 3476 4180 3572 4220
rect 3436 4171 3476 4180
rect 3532 3641 3572 4180
rect 3628 3977 3668 5104
rect 3627 3968 3669 3977
rect 3627 3928 3628 3968
rect 3668 3928 3669 3968
rect 3627 3919 3669 3928
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3531 3632 3573 3641
rect 4108 3632 4148 5440
rect 4204 4061 4244 5524
rect 4299 5524 4300 5564
rect 4340 5524 4341 5564
rect 4299 5515 4341 5524
rect 4203 4052 4245 4061
rect 4203 4012 4204 4052
rect 4244 4012 4245 4052
rect 4203 4003 4245 4012
rect 4203 3884 4245 3893
rect 4203 3844 4204 3884
rect 4244 3844 4245 3884
rect 4203 3835 4245 3844
rect 3531 3592 3532 3632
rect 3572 3592 3573 3632
rect 3531 3583 3573 3592
rect 4012 3592 4148 3632
rect 3147 3464 3189 3473
rect 3147 3424 3148 3464
rect 3188 3424 3189 3464
rect 3147 3415 3189 3424
rect 2956 3331 2996 3340
rect 3148 3380 3188 3415
rect 3148 3329 3188 3340
rect 3819 3380 3861 3389
rect 3819 3340 3820 3380
rect 3860 3340 3861 3380
rect 3819 3331 3861 3340
rect 4012 3380 4052 3592
rect 4012 3331 4052 3340
rect 4108 3380 4148 3391
rect 1899 3296 1941 3305
rect 1899 3256 1900 3296
rect 1940 3256 1941 3296
rect 1899 3247 1941 3256
rect 2571 3296 2613 3305
rect 2571 3256 2572 3296
rect 2612 3256 2613 3296
rect 2571 3247 2613 3256
rect 3820 3246 3860 3331
rect 4108 3305 4148 3340
rect 4204 3380 4244 3835
rect 4300 3389 4340 5515
rect 4588 4229 4628 5599
rect 4684 4724 4724 4733
rect 4587 4220 4629 4229
rect 4587 4180 4588 4220
rect 4628 4180 4629 4220
rect 4587 4171 4629 4180
rect 4684 4061 4724 4684
rect 4780 4397 4820 5683
rect 4972 5480 5012 5489
rect 4972 5069 5012 5440
rect 4971 5060 5013 5069
rect 4971 5020 4972 5060
rect 5012 5020 5013 5060
rect 4971 5011 5013 5020
rect 4971 4892 5013 4901
rect 4971 4852 4972 4892
rect 5012 4852 5013 4892
rect 4971 4843 5013 4852
rect 4972 4758 5012 4843
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4779 4388 4821 4397
rect 4779 4348 4780 4388
rect 4820 4348 4821 4388
rect 4779 4339 4821 4348
rect 4876 4388 4916 4397
rect 5452 4388 5492 5692
rect 5644 5683 5684 5692
rect 6027 5732 6069 5741
rect 6027 5692 6028 5732
rect 6068 5692 6069 5732
rect 6027 5683 6069 5692
rect 5547 5564 5589 5573
rect 5547 5524 5548 5564
rect 5588 5524 5589 5564
rect 5547 5515 5589 5524
rect 4876 4229 4916 4348
rect 4972 4348 5492 4388
rect 4875 4220 4917 4229
rect 4875 4180 4876 4220
rect 4916 4180 4917 4220
rect 4875 4171 4917 4180
rect 4683 4052 4725 4061
rect 4683 4012 4684 4052
rect 4724 4012 4725 4052
rect 4683 4003 4725 4012
rect 4588 3968 4628 3977
rect 4492 3557 4532 3642
rect 4491 3548 4533 3557
rect 4491 3508 4492 3548
rect 4532 3508 4533 3548
rect 4491 3499 4533 3508
rect 4588 3473 4628 3928
rect 4972 3632 5012 4348
rect 5067 4220 5109 4229
rect 5067 4180 5068 4220
rect 5108 4180 5109 4220
rect 5067 4171 5109 4180
rect 5164 4220 5204 4231
rect 5068 4086 5108 4171
rect 5164 4145 5204 4180
rect 5259 4220 5301 4229
rect 5259 4180 5260 4220
rect 5300 4180 5301 4220
rect 5259 4171 5301 4180
rect 5356 4220 5396 4229
rect 5163 4136 5205 4145
rect 5163 4096 5164 4136
rect 5204 4096 5205 4136
rect 5163 4087 5205 4096
rect 5164 3632 5204 4087
rect 5260 3977 5300 4171
rect 5259 3968 5301 3977
rect 5259 3928 5260 3968
rect 5300 3928 5301 3968
rect 5259 3919 5301 3928
rect 4972 3583 5012 3592
rect 5068 3592 5204 3632
rect 4587 3464 4629 3473
rect 4587 3424 4588 3464
rect 4628 3424 4629 3464
rect 4587 3415 4629 3424
rect 4204 3331 4244 3340
rect 4299 3380 4341 3389
rect 4299 3340 4300 3380
rect 4340 3340 4341 3380
rect 4299 3331 4341 3340
rect 4491 3380 4533 3389
rect 4491 3340 4492 3380
rect 4532 3340 4533 3380
rect 4491 3331 4533 3340
rect 4684 3380 4724 3389
rect 4107 3296 4149 3305
rect 4107 3256 4108 3296
rect 4148 3256 4149 3296
rect 4107 3247 4149 3256
rect 4300 3246 4340 3331
rect 4492 3246 4532 3331
rect 2188 3212 2228 3221
rect 4684 3212 4724 3340
rect 4780 3380 4820 3389
rect 4972 3380 5012 3389
rect 5068 3380 5108 3592
rect 5356 3557 5396 4180
rect 5355 3548 5397 3557
rect 5355 3508 5356 3548
rect 5396 3508 5397 3548
rect 5355 3499 5397 3508
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 4820 3340 4972 3380
rect 5012 3340 5108 3380
rect 5164 3380 5204 3415
rect 4780 3331 4820 3340
rect 4972 3331 5012 3340
rect 5164 3329 5204 3340
rect 5260 3380 5300 3389
rect 5548 3380 5588 5515
rect 5739 5480 5781 5489
rect 5739 5440 5740 5480
rect 5780 5440 5781 5480
rect 5739 5431 5781 5440
rect 5836 5480 5876 5489
rect 5876 5440 5972 5480
rect 5836 5431 5876 5440
rect 5740 4892 5780 5431
rect 5836 4892 5876 4901
rect 5740 4852 5836 4892
rect 5836 4843 5876 4852
rect 5644 4724 5684 4733
rect 5644 4313 5684 4684
rect 5835 4724 5877 4733
rect 5835 4684 5836 4724
rect 5876 4684 5877 4724
rect 5835 4675 5877 4684
rect 5643 4304 5685 4313
rect 5643 4264 5644 4304
rect 5684 4264 5685 4304
rect 5643 4255 5685 4264
rect 5836 4136 5876 4675
rect 5932 4229 5972 5440
rect 6028 4733 6068 5683
rect 6220 4892 6260 6103
rect 6508 5732 6548 8371
rect 7084 7916 7124 8539
rect 7084 7244 7124 7876
rect 7084 7195 7124 7204
rect 7276 6833 7316 9388
rect 7468 9379 7508 9388
rect 7468 8756 7508 8765
rect 7852 8756 7892 9472
rect 8044 9260 8084 9269
rect 8427 9260 8469 9269
rect 8084 9220 8180 9260
rect 8044 9211 8084 9220
rect 7508 8716 7892 8756
rect 7468 7421 7508 8716
rect 7660 8588 7700 8597
rect 8044 8588 8084 8597
rect 7660 7925 7700 8548
rect 7948 8548 8044 8588
rect 7659 7916 7701 7925
rect 7659 7876 7660 7916
rect 7700 7876 7701 7916
rect 7659 7867 7701 7876
rect 7467 7412 7509 7421
rect 7467 7372 7468 7412
rect 7508 7372 7509 7412
rect 7467 7363 7509 7372
rect 7948 7253 7988 8548
rect 8044 8539 8084 8548
rect 8140 8009 8180 9220
rect 8427 9220 8428 9260
rect 8468 9220 8469 9260
rect 8427 9211 8469 9220
rect 8331 8168 8373 8177
rect 8331 8128 8332 8168
rect 8372 8128 8373 8168
rect 8331 8119 8373 8128
rect 8139 8000 8181 8009
rect 8139 7960 8140 8000
rect 8180 7960 8181 8000
rect 8139 7951 8181 7960
rect 8236 7748 8276 7757
rect 8044 7708 8236 7748
rect 7947 7244 7989 7253
rect 7947 7204 7948 7244
rect 7988 7204 7989 7244
rect 7947 7195 7989 7204
rect 7275 6824 7317 6833
rect 7275 6784 7276 6824
rect 7316 6784 7317 6824
rect 7275 6775 7317 6784
rect 7179 6656 7221 6665
rect 7179 6616 7180 6656
rect 7220 6616 7221 6656
rect 7179 6607 7221 6616
rect 7180 6488 7220 6607
rect 6508 5573 6548 5692
rect 7084 6448 7220 6488
rect 8044 6488 8084 7708
rect 8236 7699 8276 7708
rect 8235 7412 8277 7421
rect 8235 7372 8236 7412
rect 8276 7372 8277 7412
rect 8235 7363 8277 7372
rect 8236 7278 8276 7363
rect 8236 6656 8276 6665
rect 8332 6656 8372 8119
rect 8276 6616 8372 6656
rect 8236 6607 8276 6616
rect 6507 5564 6549 5573
rect 6507 5524 6508 5564
rect 6548 5524 6549 5564
rect 6507 5515 6549 5524
rect 6508 5153 6548 5515
rect 6700 5480 6740 5489
rect 6507 5144 6549 5153
rect 6507 5104 6508 5144
rect 6548 5104 6549 5144
rect 6507 5095 6549 5104
rect 6220 4843 6260 4852
rect 6027 4724 6069 4733
rect 6027 4684 6028 4724
rect 6068 4684 6069 4724
rect 6027 4675 6069 4684
rect 6700 4397 6740 5440
rect 7084 5312 7124 6448
rect 7468 6404 7508 6413
rect 7852 6404 7892 6413
rect 7508 6364 7700 6404
rect 7468 6355 7508 6364
rect 7371 5732 7413 5741
rect 7371 5692 7372 5732
rect 7412 5692 7413 5732
rect 7660 5732 7700 6364
rect 7892 6364 7988 6404
rect 7852 6355 7892 6364
rect 7756 6245 7796 6330
rect 7755 6236 7797 6245
rect 7755 6196 7756 6236
rect 7796 6196 7797 6236
rect 7755 6187 7797 6196
rect 7660 5692 7796 5732
rect 7371 5683 7413 5692
rect 7372 5598 7412 5683
rect 7564 5489 7604 5574
rect 7563 5480 7605 5489
rect 7563 5440 7564 5480
rect 7604 5440 7605 5480
rect 7563 5431 7605 5440
rect 7084 5272 7508 5312
rect 7084 4892 7124 4901
rect 6699 4388 6741 4397
rect 6699 4348 6700 4388
rect 6740 4348 6741 4388
rect 6699 4339 6741 4348
rect 5931 4220 5973 4229
rect 5931 4180 5932 4220
rect 5972 4180 5973 4220
rect 5931 4171 5973 4180
rect 6988 4220 7028 4229
rect 7084 4220 7124 4852
rect 7028 4180 7124 4220
rect 5836 4087 5876 4096
rect 6988 3641 7028 4180
rect 5739 3632 5781 3641
rect 5739 3592 5740 3632
rect 5780 3592 5781 3632
rect 5739 3583 5781 3592
rect 6987 3632 7029 3641
rect 6987 3592 6988 3632
rect 7028 3592 7029 3632
rect 6987 3583 7029 3592
rect 5740 3498 5780 3583
rect 5300 3340 5588 3380
rect 7468 3380 7508 5272
rect 7756 4985 7796 5692
rect 7948 5489 7988 6364
rect 8044 5732 8084 6448
rect 8236 5732 8276 5741
rect 8044 5692 8236 5732
rect 8236 5683 8276 5692
rect 7947 5480 7989 5489
rect 7947 5440 7948 5480
rect 7988 5440 7989 5480
rect 7947 5431 7989 5440
rect 8235 5144 8277 5153
rect 8235 5104 8236 5144
rect 8276 5104 8277 5144
rect 8235 5095 8277 5104
rect 8236 5010 8276 5095
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 8428 4817 8468 9211
rect 8427 4808 8469 4817
rect 8427 4768 8428 4808
rect 8468 4768 8469 4808
rect 8427 4759 8469 4768
rect 8235 4304 8277 4313
rect 8235 4264 8236 4304
rect 8276 4264 8277 4304
rect 8235 4255 8277 4264
rect 7852 4220 7892 4229
rect 7852 3548 7892 4180
rect 8236 4170 8276 4255
rect 7852 3499 7892 3508
rect 5260 3212 5300 3340
rect 7468 3331 7508 3340
rect 4684 3172 5300 3212
rect 2188 2969 2228 3172
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 2187 2960 2229 2969
rect 2187 2920 2188 2960
rect 2228 2920 2229 2960
rect 2187 2911 2229 2920
rect 4491 2960 4533 2969
rect 4491 2920 4492 2960
rect 4532 2920 4533 2960
rect 4491 2911 4533 2920
rect 4492 80 4532 2911
rect 4472 0 4552 80
<< via2 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 1420 9472 1460 9512
rect 2476 9472 2516 9512
rect 1804 9220 1844 9260
rect 1516 8548 1556 8588
rect 1228 7960 1268 8000
rect 1228 7792 1268 7832
rect 1420 7120 1460 7160
rect 1612 7624 1652 7664
rect 1900 8716 1940 8756
rect 2380 9220 2420 9260
rect 2476 8884 2516 8924
rect 2380 8716 2420 8756
rect 2092 8044 2132 8084
rect 1804 6700 1844 6740
rect 1612 6448 1652 6488
rect 1708 6280 1748 6320
rect 1228 5692 1268 5732
rect 1708 5692 1748 5732
rect 1324 4936 1364 4976
rect 1420 4852 1460 4892
rect 1228 4516 1268 4556
rect 1708 5020 1748 5060
rect 2092 6364 2132 6404
rect 1996 6280 2036 6320
rect 1900 6196 1940 6236
rect 4012 9388 4052 9428
rect 3916 9304 3956 9344
rect 3532 8884 3572 8924
rect 3724 8884 3764 8924
rect 2668 8716 2708 8756
rect 4012 8800 4052 8840
rect 2668 8044 2708 8084
rect 3724 8716 3764 8756
rect 3916 8716 3956 8756
rect 2860 8548 2900 8588
rect 3532 8548 3572 8588
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3340 6448 3380 6488
rect 4684 9304 4724 9344
rect 4876 9388 4916 9428
rect 5260 9220 5300 9260
rect 4780 9136 4820 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4588 8884 4628 8924
rect 4780 8884 4820 8924
rect 4300 7540 4340 7580
rect 4684 8716 4724 8756
rect 6796 9136 6836 9176
rect 6604 8884 6644 8924
rect 5740 8632 5780 8672
rect 7084 8548 7124 8588
rect 5356 8380 5396 8420
rect 4492 7960 4532 8000
rect 5068 7960 5108 8000
rect 4396 7456 4436 7496
rect 4684 7456 4724 7496
rect 6508 8380 6548 8420
rect 6220 7876 6260 7916
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5164 7372 5204 7412
rect 4108 6364 4148 6404
rect 3532 6196 3572 6236
rect 2476 6112 2516 6152
rect 2380 5776 2420 5816
rect 1996 5692 2036 5732
rect 1996 5524 2036 5564
rect 1804 4936 1844 4976
rect 1612 4600 1652 4640
rect 1612 4264 1652 4304
rect 1420 3424 1460 3464
rect 1708 3340 1748 3380
rect 4588 7120 4628 7160
rect 4684 7036 4724 7076
rect 4588 6364 4628 6404
rect 4972 6448 5012 6488
rect 6220 7204 6260 7244
rect 5548 6448 5588 6488
rect 6028 6448 6068 6488
rect 5164 6364 5204 6404
rect 6220 6112 6260 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4204 5776 4244 5816
rect 2476 5692 2516 5732
rect 3340 5524 3380 5564
rect 3724 5524 3764 5564
rect 3916 5440 3956 5480
rect 4780 5692 4820 5732
rect 4588 5608 4628 5648
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 2668 5020 2708 5060
rect 2956 5020 2996 5060
rect 2764 4852 2804 4892
rect 2188 4264 2228 4304
rect 2092 4180 2132 4220
rect 1996 4012 2036 4052
rect 2572 4180 2612 4220
rect 2380 3508 2420 3548
rect 3628 3928 3668 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4300 5524 4340 5564
rect 4204 4012 4244 4052
rect 4204 3844 4244 3884
rect 3532 3592 3572 3632
rect 3148 3424 3188 3464
rect 3820 3340 3860 3380
rect 1900 3256 1940 3296
rect 2572 3256 2612 3296
rect 4588 4180 4628 4220
rect 4972 5020 5012 5060
rect 4972 4852 5012 4892
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4780 4348 4820 4388
rect 6028 5692 6068 5732
rect 5548 5524 5588 5564
rect 4876 4180 4916 4220
rect 4684 4012 4724 4052
rect 4492 3508 4532 3548
rect 5068 4180 5108 4220
rect 5260 4180 5300 4220
rect 5164 4096 5204 4136
rect 5260 3928 5300 3968
rect 4588 3424 4628 3464
rect 4300 3340 4340 3380
rect 4492 3340 4532 3380
rect 4108 3256 4148 3296
rect 5356 3508 5396 3548
rect 5164 3424 5204 3464
rect 5740 5440 5780 5480
rect 5836 4684 5876 4724
rect 5644 4264 5684 4304
rect 7660 7876 7700 7916
rect 7468 7372 7508 7412
rect 8428 9220 8468 9260
rect 8332 8128 8372 8168
rect 8140 7960 8180 8000
rect 7948 7204 7988 7244
rect 7276 6784 7316 6824
rect 7180 6616 7220 6656
rect 8236 7372 8276 7412
rect 6508 5524 6548 5564
rect 6508 5104 6548 5144
rect 6028 4684 6068 4724
rect 7372 5692 7412 5732
rect 7756 6196 7796 6236
rect 7564 5440 7604 5480
rect 6700 4348 6740 4388
rect 5932 4180 5972 4220
rect 5740 3592 5780 3632
rect 6988 3592 7028 3632
rect 7948 5440 7988 5480
rect 8236 5104 8276 5144
rect 7756 4936 7796 4976
rect 8428 4768 8468 4808
rect 8236 4264 8276 4304
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 2188 2920 2228 2960
rect 4492 2920 4532 2960
<< metal3 >>
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 1411 9472 1420 9512
rect 1460 9472 2476 9512
rect 2516 9472 2525 9512
rect 4003 9388 4012 9428
rect 4052 9388 4876 9428
rect 4916 9388 4925 9428
rect 3907 9304 3916 9344
rect 3956 9304 4684 9344
rect 4724 9304 4733 9344
rect 1795 9220 1804 9260
rect 1844 9220 2380 9260
rect 2420 9220 2429 9260
rect 5251 9220 5260 9260
rect 5300 9220 8428 9260
rect 8468 9220 8477 9260
rect 4675 9176 4733 9177
rect 4675 9136 4684 9176
rect 4724 9136 4780 9176
rect 4820 9136 6796 9176
rect 6836 9136 6845 9176
rect 4675 9135 4733 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 4579 8924 4637 8925
rect 2467 8884 2476 8924
rect 2516 8884 3532 8924
rect 3572 8884 3724 8924
rect 3764 8884 4588 8924
rect 4628 8884 4637 8924
rect 4771 8884 4780 8924
rect 4820 8884 6604 8924
rect 6644 8884 6653 8924
rect 4579 8883 4637 8884
rect 2380 8800 4012 8840
rect 4052 8800 4061 8840
rect 2380 8756 2420 8800
rect 4771 8756 4829 8757
rect 1891 8716 1900 8756
rect 1940 8716 2380 8756
rect 2420 8716 2429 8756
rect 2659 8716 2668 8756
rect 2708 8716 3724 8756
rect 3764 8716 3916 8756
rect 3956 8716 3965 8756
rect 4675 8716 4684 8756
rect 4724 8716 4780 8756
rect 4820 8716 4829 8756
rect 4771 8715 4829 8716
rect 5731 8632 5740 8672
rect 5780 8632 5789 8672
rect 5740 8588 5780 8632
rect 1507 8548 1516 8588
rect 1556 8548 2860 8588
rect 2900 8548 2909 8588
rect 3523 8548 3532 8588
rect 3572 8548 7084 8588
rect 7124 8548 7133 8588
rect 5347 8380 5356 8420
rect 5396 8380 6508 8420
rect 6548 8380 6557 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 9483 8168 9563 8188
rect 8323 8128 8332 8168
rect 8372 8128 9563 8168
rect 9483 8108 9563 8128
rect 2083 8044 2092 8084
rect 2132 8044 2668 8084
rect 2708 8044 2717 8084
rect 0 8000 80 8020
rect 9483 8000 9563 8020
rect 0 7960 1228 8000
rect 1268 7960 1277 8000
rect 4483 7960 4492 8000
rect 4532 7960 5068 8000
rect 5108 7960 5117 8000
rect 8131 7960 8140 8000
rect 8180 7960 9563 8000
rect 0 7940 80 7960
rect 9483 7940 9563 7960
rect 6211 7876 6220 7916
rect 6260 7876 7660 7916
rect 7700 7876 7709 7916
rect 0 7832 80 7852
rect 0 7792 1228 7832
rect 1268 7792 1277 7832
rect 0 7772 80 7792
rect 0 7664 80 7684
rect 0 7624 1612 7664
rect 1652 7624 1661 7664
rect 0 7604 80 7624
rect 4291 7540 4300 7580
rect 4340 7540 4820 7580
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 4301 7456 4396 7496
rect 4436 7456 4684 7496
rect 4724 7456 4733 7496
rect 4396 7160 4436 7456
rect 4780 7412 4820 7540
rect 4780 7372 5164 7412
rect 5204 7372 5213 7412
rect 7459 7372 7468 7412
rect 7508 7372 8236 7412
rect 8276 7372 8285 7412
rect 6211 7204 6220 7244
rect 6260 7204 7948 7244
rect 7988 7204 7997 7244
rect 1411 7120 1420 7160
rect 1460 7120 4436 7160
rect 4579 7160 4637 7161
rect 4579 7120 4588 7160
rect 4628 7120 4722 7160
rect 4579 7119 4637 7120
rect 4675 7076 4733 7077
rect 4590 7036 4684 7076
rect 4724 7036 4733 7076
rect 4675 7035 4733 7036
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 7180 6784 7276 6824
rect 7316 6784 7325 6824
rect 1795 6700 1804 6740
rect 1844 6700 2900 6740
rect 2860 6572 2900 6700
rect 7180 6656 7220 6784
rect 7171 6616 7180 6656
rect 7220 6616 7315 6656
rect 2860 6532 5012 6572
rect 4972 6488 5012 6532
rect 7180 6488 7220 6616
rect 1603 6448 1612 6488
rect 1652 6448 3340 6488
rect 3380 6448 3389 6488
rect 4963 6448 4972 6488
rect 5012 6448 5548 6488
rect 5588 6448 5597 6488
rect 6019 6448 6028 6488
rect 6068 6448 7220 6488
rect 4771 6404 4829 6405
rect 2083 6364 2092 6404
rect 2132 6364 4108 6404
rect 4148 6364 4588 6404
rect 4628 6364 4637 6404
rect 4771 6364 4780 6404
rect 4820 6364 5164 6404
rect 5204 6364 5213 6404
rect 4771 6363 4829 6364
rect 1699 6280 1708 6320
rect 1748 6280 1996 6320
rect 2036 6280 2045 6320
rect 5164 6236 5204 6364
rect 1891 6196 1900 6236
rect 1940 6196 3532 6236
rect 3572 6196 3581 6236
rect 5164 6196 7756 6236
rect 7796 6196 7805 6236
rect 2467 6112 2476 6152
rect 2516 6112 6220 6152
rect 6260 6112 6269 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 2371 5776 2380 5816
rect 2420 5776 4204 5816
rect 4244 5776 4253 5816
rect 1219 5692 1228 5732
rect 1268 5692 1708 5732
rect 1748 5692 1757 5732
rect 1987 5692 1996 5732
rect 2036 5692 2045 5732
rect 2467 5692 2476 5732
rect 2516 5692 4780 5732
rect 4820 5692 4829 5732
rect 6019 5692 6028 5732
rect 6068 5692 7372 5732
rect 7412 5692 7421 5732
rect 1996 5648 2036 5692
rect 1996 5608 4588 5648
rect 4628 5608 4637 5648
rect 1987 5524 1996 5564
rect 2036 5524 3340 5564
rect 3380 5524 3389 5564
rect 3715 5524 3724 5564
rect 3764 5524 4300 5564
rect 4340 5524 4349 5564
rect 5539 5524 5548 5564
rect 5588 5524 6508 5564
rect 6548 5524 6557 5564
rect 3907 5440 3916 5480
rect 3956 5440 5740 5480
rect 5780 5440 5789 5480
rect 7555 5440 7564 5480
rect 7604 5440 7948 5480
rect 7988 5440 7997 5480
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 6499 5104 6508 5144
rect 6548 5104 8236 5144
rect 8276 5104 8285 5144
rect 1699 5020 1708 5060
rect 1748 5020 2668 5060
rect 2708 5020 2717 5060
rect 2947 5020 2956 5060
rect 2996 5020 4972 5060
rect 5012 5020 5021 5060
rect 9483 4976 9563 4996
rect 1315 4936 1324 4976
rect 1364 4936 1804 4976
rect 1844 4936 1853 4976
rect 7747 4936 7756 4976
rect 7796 4936 9563 4976
rect 9483 4916 9563 4936
rect 1411 4852 1420 4892
rect 1460 4852 1469 4892
rect 2755 4852 2764 4892
rect 2804 4852 4972 4892
rect 5012 4852 5021 4892
rect 1420 4724 1460 4852
rect 9483 4808 9563 4828
rect 8419 4768 8428 4808
rect 8468 4768 9563 4808
rect 9483 4748 9563 4768
rect 1420 4684 5836 4724
rect 5876 4684 6028 4724
rect 6068 4684 6077 4724
rect 0 4640 80 4660
rect 9483 4640 9563 4660
rect 0 4600 1268 4640
rect 1603 4600 1612 4640
rect 1652 4600 9563 4640
rect 0 4580 80 4600
rect 1228 4556 1268 4600
rect 9483 4580 9563 4600
rect 1219 4516 1228 4556
rect 1268 4516 1277 4556
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 4771 4348 4780 4388
rect 4820 4348 5108 4388
rect 1603 4264 1612 4304
rect 1652 4264 2188 4304
rect 2228 4264 2237 4304
rect 5068 4220 5108 4348
rect 5164 4348 6700 4388
rect 6740 4348 6749 4388
rect 2083 4180 2092 4220
rect 2132 4180 2572 4220
rect 2612 4180 2621 4220
rect 4579 4180 4588 4220
rect 4628 4180 4876 4220
rect 4916 4180 4925 4220
rect 5059 4180 5068 4220
rect 5108 4180 5117 4220
rect 5164 4136 5204 4348
rect 5635 4264 5644 4304
rect 5684 4264 8236 4304
rect 8276 4264 8285 4304
rect 5251 4180 5260 4220
rect 5300 4180 5932 4220
rect 5972 4180 5981 4220
rect 5155 4096 5164 4136
rect 5204 4096 5213 4136
rect 1987 4012 1996 4052
rect 2036 4012 4204 4052
rect 4244 4012 4684 4052
rect 4724 4012 4733 4052
rect 3619 3928 3628 3968
rect 3668 3928 5260 3968
rect 5300 3928 5309 3968
rect 4204 3884 4244 3928
rect 4195 3844 4204 3884
rect 4244 3844 4284 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 3523 3592 3532 3632
rect 3572 3592 5740 3632
rect 5780 3592 6988 3632
rect 7028 3592 7037 3632
rect 2371 3508 2380 3548
rect 2420 3508 4492 3548
rect 4532 3508 4541 3548
rect 5347 3508 5356 3548
rect 5396 3508 5405 3548
rect 1411 3424 1420 3464
rect 1460 3424 3148 3464
rect 3188 3424 4588 3464
rect 4628 3424 5164 3464
rect 5204 3424 5213 3464
rect 5356 3380 5396 3508
rect 1699 3340 1708 3380
rect 1748 3340 3820 3380
rect 3860 3340 4300 3380
rect 4340 3340 4492 3380
rect 4532 3340 5396 3380
rect 1891 3256 1900 3296
rect 1940 3256 2572 3296
rect 2612 3256 4108 3296
rect 4148 3256 4157 3296
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 2179 2920 2188 2960
rect 2228 2920 4492 2960
rect 4532 2920 4541 2960
<< via3 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4684 9136 4724 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4588 8884 4628 8924
rect 4780 8716 4820 8756
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4588 7120 4628 7160
rect 4684 7036 4724 7076
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4780 6364 4820 6404
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal4 >>
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4684 9176 4724 9185
rect 4588 8924 4628 8933
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4588 7160 4628 8884
rect 4588 7111 4628 7120
rect 4684 7076 4724 9136
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4684 7027 4724 7036
rect 4780 8756 4820 8765
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4780 6404 4820 8716
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4780 6355 4820 6364
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
<< metal5 >>
rect 3679 9848 3726 9890
rect 3850 9848 3894 9890
rect 4018 9848 4065 9890
rect 3679 9808 3688 9848
rect 3850 9808 3852 9848
rect 3892 9808 3894 9848
rect 4056 9808 4065 9848
rect 3679 9766 3726 9808
rect 3850 9766 3894 9808
rect 4018 9766 4065 9808
rect 4919 9092 4966 9134
rect 5090 9092 5134 9134
rect 5258 9092 5305 9134
rect 4919 9052 4928 9092
rect 5090 9052 5092 9092
rect 5132 9052 5134 9092
rect 5296 9052 5305 9092
rect 4919 9010 4966 9052
rect 5090 9010 5134 9052
rect 5258 9010 5305 9052
rect 3679 8336 3726 8378
rect 3850 8336 3894 8378
rect 4018 8336 4065 8378
rect 3679 8296 3688 8336
rect 3850 8296 3852 8336
rect 3892 8296 3894 8336
rect 4056 8296 4065 8336
rect 3679 8254 3726 8296
rect 3850 8254 3894 8296
rect 4018 8254 4065 8296
rect 4919 7580 4966 7622
rect 5090 7580 5134 7622
rect 5258 7580 5305 7622
rect 4919 7540 4928 7580
rect 5090 7540 5092 7580
rect 5132 7540 5134 7580
rect 5296 7540 5305 7580
rect 4919 7498 4966 7540
rect 5090 7498 5134 7540
rect 5258 7498 5305 7540
rect 3679 6824 3726 6866
rect 3850 6824 3894 6866
rect 4018 6824 4065 6866
rect 3679 6784 3688 6824
rect 3850 6784 3852 6824
rect 3892 6784 3894 6824
rect 4056 6784 4065 6824
rect 3679 6742 3726 6784
rect 3850 6742 3894 6784
rect 4018 6742 4065 6784
rect 4919 6068 4966 6110
rect 5090 6068 5134 6110
rect 5258 6068 5305 6110
rect 4919 6028 4928 6068
rect 5090 6028 5092 6068
rect 5132 6028 5134 6068
rect 5296 6028 5305 6068
rect 4919 5986 4966 6028
rect 5090 5986 5134 6028
rect 5258 5986 5305 6028
rect 3679 5312 3726 5354
rect 3850 5312 3894 5354
rect 4018 5312 4065 5354
rect 3679 5272 3688 5312
rect 3850 5272 3852 5312
rect 3892 5272 3894 5312
rect 4056 5272 4065 5312
rect 3679 5230 3726 5272
rect 3850 5230 3894 5272
rect 4018 5230 4065 5272
rect 4919 4556 4966 4598
rect 5090 4556 5134 4598
rect 5258 4556 5305 4598
rect 4919 4516 4928 4556
rect 5090 4516 5092 4556
rect 5132 4516 5134 4556
rect 5296 4516 5305 4556
rect 4919 4474 4966 4516
rect 5090 4474 5134 4516
rect 5258 4474 5305 4516
rect 3679 3800 3726 3842
rect 3850 3800 3894 3842
rect 4018 3800 4065 3842
rect 3679 3760 3688 3800
rect 3850 3760 3852 3800
rect 3892 3760 3894 3800
rect 4056 3760 4065 3800
rect 3679 3718 3726 3760
rect 3850 3718 3894 3760
rect 4018 3718 4065 3760
rect 4919 3044 4966 3086
rect 5090 3044 5134 3086
rect 5258 3044 5305 3086
rect 4919 3004 4928 3044
rect 5090 3004 5092 3044
rect 5132 3004 5134 3044
rect 5296 3004 5305 3044
rect 4919 2962 4966 3004
rect 5090 2962 5134 3004
rect 5258 2962 5305 3004
<< via5 >>
rect 3726 9848 3850 9890
rect 3894 9848 4018 9890
rect 3726 9808 3728 9848
rect 3728 9808 3770 9848
rect 3770 9808 3810 9848
rect 3810 9808 3850 9848
rect 3894 9808 3934 9848
rect 3934 9808 3974 9848
rect 3974 9808 4016 9848
rect 4016 9808 4018 9848
rect 3726 9766 3850 9808
rect 3894 9766 4018 9808
rect 4966 9092 5090 9134
rect 5134 9092 5258 9134
rect 4966 9052 4968 9092
rect 4968 9052 5010 9092
rect 5010 9052 5050 9092
rect 5050 9052 5090 9092
rect 5134 9052 5174 9092
rect 5174 9052 5214 9092
rect 5214 9052 5256 9092
rect 5256 9052 5258 9092
rect 4966 9010 5090 9052
rect 5134 9010 5258 9052
rect 3726 8336 3850 8378
rect 3894 8336 4018 8378
rect 3726 8296 3728 8336
rect 3728 8296 3770 8336
rect 3770 8296 3810 8336
rect 3810 8296 3850 8336
rect 3894 8296 3934 8336
rect 3934 8296 3974 8336
rect 3974 8296 4016 8336
rect 4016 8296 4018 8336
rect 3726 8254 3850 8296
rect 3894 8254 4018 8296
rect 4966 7580 5090 7622
rect 5134 7580 5258 7622
rect 4966 7540 4968 7580
rect 4968 7540 5010 7580
rect 5010 7540 5050 7580
rect 5050 7540 5090 7580
rect 5134 7540 5174 7580
rect 5174 7540 5214 7580
rect 5214 7540 5256 7580
rect 5256 7540 5258 7580
rect 4966 7498 5090 7540
rect 5134 7498 5258 7540
rect 3726 6824 3850 6866
rect 3894 6824 4018 6866
rect 3726 6784 3728 6824
rect 3728 6784 3770 6824
rect 3770 6784 3810 6824
rect 3810 6784 3850 6824
rect 3894 6784 3934 6824
rect 3934 6784 3974 6824
rect 3974 6784 4016 6824
rect 4016 6784 4018 6824
rect 3726 6742 3850 6784
rect 3894 6742 4018 6784
rect 4966 6068 5090 6110
rect 5134 6068 5258 6110
rect 4966 6028 4968 6068
rect 4968 6028 5010 6068
rect 5010 6028 5050 6068
rect 5050 6028 5090 6068
rect 5134 6028 5174 6068
rect 5174 6028 5214 6068
rect 5214 6028 5256 6068
rect 5256 6028 5258 6068
rect 4966 5986 5090 6028
rect 5134 5986 5258 6028
rect 3726 5312 3850 5354
rect 3894 5312 4018 5354
rect 3726 5272 3728 5312
rect 3728 5272 3770 5312
rect 3770 5272 3810 5312
rect 3810 5272 3850 5312
rect 3894 5272 3934 5312
rect 3934 5272 3974 5312
rect 3974 5272 4016 5312
rect 4016 5272 4018 5312
rect 3726 5230 3850 5272
rect 3894 5230 4018 5272
rect 4966 4556 5090 4598
rect 5134 4556 5258 4598
rect 4966 4516 4968 4556
rect 4968 4516 5010 4556
rect 5010 4516 5050 4556
rect 5050 4516 5090 4556
rect 5134 4516 5174 4556
rect 5174 4516 5214 4556
rect 5214 4516 5256 4556
rect 5256 4516 5258 4556
rect 4966 4474 5090 4516
rect 5134 4474 5258 4516
rect 3726 3800 3850 3842
rect 3894 3800 4018 3842
rect 3726 3760 3728 3800
rect 3728 3760 3770 3800
rect 3770 3760 3810 3800
rect 3810 3760 3850 3800
rect 3894 3760 3934 3800
rect 3934 3760 3974 3800
rect 3974 3760 4016 3800
rect 4016 3760 4018 3800
rect 3726 3718 3850 3760
rect 3894 3718 4018 3760
rect 4966 3044 5090 3086
rect 5134 3044 5258 3086
rect 4966 3004 4968 3044
rect 4968 3004 5010 3044
rect 5010 3004 5050 3044
rect 5050 3004 5090 3044
rect 5134 3004 5174 3044
rect 5174 3004 5214 3044
rect 5214 3004 5256 3044
rect 5256 3004 5258 3044
rect 4966 2962 5090 3004
rect 5134 2962 5258 3004
<< metal6 >>
rect 3652 9890 4092 9954
rect 3652 9766 3726 9890
rect 3850 9766 3894 9890
rect 4018 9766 4092 9890
rect 3652 8378 4092 9766
rect 3652 8254 3726 8378
rect 3850 8254 3894 8378
rect 4018 8254 4092 8378
rect 3652 6866 4092 8254
rect 3652 6742 3726 6866
rect 3850 6742 3894 6866
rect 4018 6742 4092 6866
rect 3652 5934 4092 6742
rect 3652 5554 3682 5934
rect 4062 5554 4092 5934
rect 3652 5354 4092 5554
rect 3652 5230 3726 5354
rect 3850 5230 3894 5354
rect 4018 5230 4092 5354
rect 3652 3842 4092 5230
rect 3652 3718 3726 3842
rect 3850 3718 3894 3842
rect 4018 3718 4092 3842
rect 3652 2980 4092 3718
rect 4892 9134 5332 9872
rect 4892 9010 4966 9134
rect 5090 9010 5134 9134
rect 5258 9010 5332 9134
rect 4892 7622 5332 9010
rect 4892 7498 4966 7622
rect 5090 7498 5134 7622
rect 5258 7498 5332 7622
rect 4892 7174 5332 7498
rect 4892 6794 4922 7174
rect 5302 6794 5332 7174
rect 4892 6110 5332 6794
rect 4892 5986 4966 6110
rect 5090 5986 5134 6110
rect 5258 5986 5332 6110
rect 4892 4598 5332 5986
rect 4892 4474 4966 4598
rect 5090 4474 5134 4598
rect 5258 4474 5332 4598
rect 4892 3086 5332 4474
rect 4892 2962 4966 3086
rect 5090 2962 5134 3086
rect 5258 2962 5332 3086
rect 4892 2898 5332 2962
<< via6 >>
rect 3682 5554 4062 5934
rect 4922 6794 5302 7174
<< metal7 >>
rect 1152 7174 8352 7204
rect 1152 6794 4922 7174
rect 5302 6794 8352 7174
rect 1152 6764 8352 6794
rect 1152 5934 8352 5964
rect 1152 5554 3682 5934
rect 4062 5554 8352 5934
rect 1152 5524 8352 5554
use sg13g2_inv_1  _31_
timestamp 1676382929
transform -1 0 7968 0 1 6048
box -48 -56 336 834
use sg13g2_inv_1  _32_
timestamp 1676382929
transform -1 0 1440 0 1 4536
box -48 -56 336 834
use sg13g2_nor2_1  _33_
timestamp 1676627187
transform -1 0 1824 0 -1 4536
box -48 -56 432 834
use sg13g2_o21ai_1  _34_
timestamp 1685175443
transform -1 0 4416 0 1 3024
box -48 -56 538 834
use sg13g2_a21oi_1  _35_
timestamp 1683973020
transform -1 0 4032 0 -1 6048
box -48 -56 528 834
use sg13g2_a21oi_1  _36_
timestamp 1683973020
transform 1 0 4896 0 1 3024
box -48 -56 528 834
use sg13g2_nand3_1  _37_
timestamp 1683988354
transform -1 0 4896 0 1 3024
box -48 -56 528 834
use sg13g2_nand2_1  _38_
timestamp 1676557249
transform 1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_nor2_1  _39_
timestamp 1676627187
transform -1 0 3072 0 1 3024
box -48 -56 432 834
use sg13g2_nor2b_1  _40_
timestamp 1685181386
transform 1 0 2112 0 -1 6048
box -54 -56 528 834
use sg13g2_and4_1  _41_
timestamp 1676985977
transform -1 0 5568 0 -1 4536
box -48 -56 816 834
use sg13g2_nor3_1  _42_
timestamp 1676639442
transform 1 0 1632 0 -1 6048
box -48 -56 528 834
use sg13g2_xor2_1  _43_
timestamp 1677577977
transform 1 0 1440 0 -1 9072
box -48 -56 816 834
use sg13g2_and2_1  _44_
timestamp 1676901763
transform -1 0 2496 0 1 9072
box -48 -56 528 834
use sg13g2_a21oi_1  _45_
timestamp 1683973020
transform -1 0 2784 0 -1 9072
box -48 -56 528 834
use sg13g2_nand3_1  _46_
timestamp 1683988354
transform -1 0 4128 0 1 9072
box -48 -56 528 834
use sg13g2_nand2_1  _47_
timestamp 1676557249
transform -1 0 2208 0 1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _48_
timestamp 1676627187
transform 1 0 1440 0 1 6048
box -48 -56 432 834
use sg13g2_nand2b_1  _49_
timestamp 1676567195
transform -1 0 4800 0 1 6048
box -48 -56 528 834
use sg13g2_nand4_1  _50_
timestamp 1685201930
transform -1 0 4992 0 1 9072
box -48 -56 624 834
use sg13g2_and3_1  _51_
timestamp 1676971669
transform -1 0 5664 0 -1 7560
box -48 -56 720 834
use sg13g2_o21ai_1  _52_
timestamp 1685175443
transform -1 0 5280 0 1 6048
box -48 -56 538 834
use sg13g2_a21oi_1  _53_
timestamp 1683973020
transform -1 0 4992 0 -1 9072
box -48 -56 528 834
use sg13g2_tiehi  _54__10
timestamp 1680000651
transform 1 0 1824 0 1 4536
box -48 -56 432 834
use sg13g2_dfrbpq_1  _54_
timestamp 1746535128
transform 1 0 2112 0 -1 4536
box -48 -56 2640 834
use sg13g2_tiehi  _55__17
timestamp 1680000651
transform 1 0 2208 0 1 6048
box -48 -56 432 834
use sg13g2_dfrbpq_1  _55_
timestamp 1746535128
transform 1 0 5760 0 1 4536
box -48 -56 2640 834
use sg13g2_tiehi  _56__16
timestamp 1680000651
transform -1 0 8160 0 1 3024
box -48 -56 432 834
use sg13g2_dfrbpq_1  _56_
timestamp 1746535128
transform -1 0 8352 0 -1 4536
box -48 -56 2640 834
use sg13g2_tiehi  _57__15
timestamp 1680000651
transform 1 0 1440 0 1 4536
box -48 -56 432 834
use sg13g2_dfrbpq_1  _57_
timestamp 1746535128
transform 1 0 2208 0 1 4536
box -48 -56 2640 834
use sg13g2_tiehi  _58__14
timestamp 1680000651
transform -1 0 2976 0 1 9072
box -48 -56 432 834
use sg13g2_dfrbpq_1  _58_
timestamp 1746535128
transform 1 0 2112 0 -1 7560
box -48 -56 2640 834
use sg13g2_tiehi  _59__13
timestamp 1680000651
transform -1 0 3360 0 1 9072
box -48 -56 432 834
use sg13g2_dfrbpq_1  _59_
timestamp 1746535128
transform 1 0 2208 0 1 7560
box -48 -56 2640 834
use sg13g2_tiehi  _60__12
timestamp 1680000651
transform -1 0 8352 0 -1 9072
box -48 -56 432 834
use sg13g2_dfrbpq_1  _60_
timestamp 1746535128
transform 1 0 5760 0 -1 7560
box -48 -56 2640 834
use sg13g2_tiehi  _61__11
timestamp 1680000651
transform -1 0 7968 0 -1 9072
box -48 -56 432 834
use sg13g2_dfrbpq_1  _61_
timestamp 1746535128
transform 1 0 5760 0 1 7560
box -48 -56 2640 834
use sg13g2_buf_16  clkbuf_0_clk_i
timestamp 1676553496
transform 1 0 5280 0 1 6048
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk_i
timestamp 1676553496
transform 1 0 5376 0 1 3024
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk_i
timestamp 1676553496
transform 1 0 5376 0 1 9072
box -48 -56 2448 834
use sg13g2_decap_4  FILLER_0_4
timestamp 1679577901
transform 1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_73
timestamp 1677580104
transform 1 0 8160 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_2
timestamp 1677579658
transform 1 0 1344 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_7
timestamp 1677580104
transform 1 0 1824 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_9
timestamp 1677579658
transform 1 0 2016 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_37
timestamp 1677579658
transform 1 0 4704 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_46
timestamp 1677580104
transform 1 0 5568 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_38
timestamp 1677579658
transform 1 0 4800 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_0
timestamp 1677579658
transform 1 0 1152 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_24
timestamp 1677579658
transform 1 0 3456 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1677580104
transform 1 0 1152 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_2
timestamp 1677579658
transform 1 0 1344 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_8
timestamp 1677580104
transform 1 0 1920 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_37
timestamp 1677580104
transform 1 0 4704 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_39
timestamp 1677579658
transform 1 0 4896 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_47
timestamp 1677579658
transform 1 0 5664 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 1152 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_38
timestamp 1677579658
transform 1 0 4800 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_0
timestamp 1677580104
transform 1 0 1152 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_2
timestamp 1677579658
transform 1 0 1344 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_11
timestamp 1677579658
transform 1 0 2208 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_4
timestamp 1679577901
transform 1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_8
timestamp 1677579658
transform 1 0 1920 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_14
timestamp 1677579658
transform 1 0 2496 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_23
timestamp 1677580104
transform 1 0 3360 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_25
timestamp 1677579658
transform 1 0 3552 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_31
timestamp 1677580104
transform 1 0 4128 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_33
timestamp 1677579658
transform 1 0 4320 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_73
timestamp 1677580104
transform 1 0 8160 0 1 9072
box -48 -56 240 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677672058
transform -1 0 8352 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677672058
transform -1 0 6720 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677672058
transform -1 0 7488 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677672058
transform -1 0 5760 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677672058
transform 1 0 4896 0 1 4536
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677672058
transform 1 0 3072 0 1 3024
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677672058
transform 1 0 4032 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677672058
transform -1 0 4320 0 1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677672058
transform -1 0 3456 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677672058
transform -1 0 4512 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677672058
transform -1 0 2208 0 1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677672058
transform -1 0 3456 0 1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677672058
transform -1 0 6624 0 -1 6048
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677672058
transform -1 0 7584 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677672058
transform 1 0 4992 0 -1 9072
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677672058
transform 1 0 4896 0 1 7560
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677672058
transform -1 0 3648 0 -1 9072
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform -1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 4992 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 1248 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 1920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform -1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 7776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 7968 0 1 6048
box -48 -56 432 834
<< labels >>
flabel metal6 s 4892 2898 5332 9872 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 1152 6764 8352 7204 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3652 2980 4092 9954 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 1152 5524 8352 5964 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 9483 4916 9563 4996 0 FreeSans 320 0 0 0 clk_i
port 2 nsew signal input
flabel metal3 s 0 4580 80 4660 0 FreeSans 320 0 0 0 count_o[0]
port 3 nsew signal output
flabel metal3 s 9483 4748 9563 4828 0 FreeSans 320 0 0 0 count_o[1]
port 4 nsew signal output
flabel metal3 s 9483 4580 9563 4660 0 FreeSans 320 0 0 0 count_o[2]
port 5 nsew signal output
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 count_o[3]
port 6 nsew signal output
flabel metal3 s 0 7940 80 8020 0 FreeSans 320 0 0 0 count_o[4]
port 7 nsew signal output
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 count_o[5]
port 8 nsew signal output
flabel metal3 s 9483 7940 9563 8020 0 FreeSans 320 0 0 0 count_o[6]
port 9 nsew signal output
flabel metal3 s 9483 8108 9563 8188 0 FreeSans 320 0 0 0 count_o[7]
port 10 nsew signal output
flabel metal3 s 0 7604 80 7684 0 FreeSans 320 0 0 0 rst_ni
port 11 nsew signal input
rlabel metal1 4752 9072 4752 9072 0 VGND
rlabel metal1 4752 9828 4752 9828 0 VPWR
rlabel metal3 1920 4284 1920 4284 0 _00_
rlabel metal2 5808 4872 5808 4872 0 _01_
rlabel metal2 2880 3528 2880 3528 0 _02_
rlabel metal2 3360 5628 3360 5628 0 _03_
rlabel metal2 2208 7770 2208 7770 0 _04_
rlabel metal2 3360 6426 3360 6426 0 _05_
rlabel metal2 5088 7350 5088 7350 0 _06_
rlabel metal2 6624 8820 6624 8820 0 _07_
rlabel metal3 4992 6384 4992 6384 0 _08_
rlabel metal2 1248 5418 1248 5418 0 _09_
rlabel metal2 4032 3486 4032 3486 0 _10_
rlabel metal2 4992 3990 4992 3990 0 _11_
rlabel metal2 2400 4032 2400 4032 0 _12_
rlabel metal2 2784 3444 2784 3444 0 _13_
rlabel metal2 4224 6090 4224 6090 0 _14_
rlabel metal2 4608 4914 4608 4914 0 _15_
rlabel metal2 2016 9156 2016 9156 0 _16_
rlabel metal2 2112 7980 2112 7980 0 _17_
rlabel metal2 4032 9576 4032 9576 0 _18_
rlabel metal2 1728 6342 1728 6342 0 _19_
rlabel metal2 4416 6708 4416 6708 0 _20_
rlabel metal2 5088 6792 5088 6792 0 _21_
rlabel metal2 4752 7308 4752 7308 0 _22_
rlabel metal3 8630 4956 8630 4956 0 clk_i
rlabel metal2 7104 5880 7104 5880 0 clknet_0_clk_i
rlabel metal2 3504 4200 3504 4200 0 clknet_1_0__leaf_clk_i
rlabel metal2 3504 7896 3504 7896 0 clknet_1_1__leaf_clk_i
rlabel metal2 1248 4074 1248 4074 0 count_o[0]
rlabel metal3 8966 4788 8966 4788 0 count_o[1]
rlabel metal2 1632 5040 1632 5040 0 count_o[2]
rlabel metal2 4512 1500 4512 1500 0 count_o[3]
rlabel metal3 654 7980 654 7980 0 count_o[4]
rlabel metal2 1248 7434 1248 7434 0 count_o[5]
rlabel metal3 8822 7980 8822 7980 0 count_o[6]
rlabel metal2 8304 6636 8304 6636 0 count_o[7]
rlabel metal2 2112 4620 2112 4620 0 net
rlabel metal2 4992 6426 4992 6426 0 net1
rlabel metal2 7680 8232 7680 8232 0 net10
rlabel metal2 7968 7896 7968 7896 0 net11
rlabel metal2 3072 9156 3072 9156 0 net12
rlabel metal2 2640 9576 2640 9576 0 net13
rlabel metal3 2208 5040 2208 5040 0 net14
rlabel metal2 7872 3864 7872 3864 0 net15
rlabel metal2 6240 5502 6240 5502 0 net16
rlabel metal3 7776 5460 7776 5460 0 net17
rlabel metal2 5904 7896 5904 7896 0 net18
rlabel metal2 5184 4158 5184 4158 0 net19
rlabel metal2 3168 3402 3168 3402 0 net2
rlabel metal2 2976 4200 2976 4200 0 net20
rlabel metal2 5664 4494 5664 4494 0 net21
rlabel metal3 4080 3360 4080 3360 0 net22
rlabel metal3 5088 4284 5088 4284 0 net23
rlabel metal2 1920 5964 1920 5964 0 net24
rlabel metal2 2448 4872 2448 4872 0 net25
rlabel metal2 3936 9072 3936 9072 0 net26
rlabel metal2 1536 7056 1536 7056 0 net27
rlabel metal2 2688 6804 2688 6804 0 net28
rlabel metal3 5616 4200 5616 4200 0 net29
rlabel metal2 5280 3276 5280 3276 0 net3
rlabel metal2 4704 6720 4704 6720 0 net30
rlabel metal2 5376 7476 5376 7476 0 net31
rlabel metal2 5856 7518 5856 7518 0 net32
rlabel metal2 1536 8652 1536 8652 0 net33
rlabel metal2 5856 4410 5856 4410 0 net4
rlabel metal2 4704 4368 4704 4368 0 net5
rlabel metal2 4608 9072 4608 9072 0 net6
rlabel metal2 4704 7602 4704 7602 0 net7
rlabel metal2 7488 8064 7488 8064 0 net8
rlabel metal2 8064 6090 8064 6090 0 net9
rlabel metal3 846 7644 846 7644 0 rst_ni
<< properties >>
string FIXED_BBOX 0 0 9563 13307
<< end >>
